// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Tue Jan 12 00:34:58 2021
//
// Verilog Description of module Master
//

module Master (CLK, UART_RX, UART_TX, Matrix_DATA_Out, Matrix_LINE_SEL_Out, 
            Matrix_CTRL_Out, SRAM_OE, SRAM_WE, SRAM_CE, SRAM_DATA, 
            SRAM_ADDR, PIC_OE, PIC_WE_IN, PIC_CS, PIC_ADDR_IN, PIC_DATA_IN, 
            PIC_READY, LED);   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(6[8:14])
    input CLK;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    input UART_RX;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(10[3:10])
    output UART_TX;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(11[3:10])
    output [11:0]Matrix_DATA_Out;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    output [3:0]Matrix_LINE_SEL_Out;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    output [2:0]Matrix_CTRL_Out;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    output SRAM_OE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(17[3:10])
    output SRAM_WE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(18[3:10])
    output SRAM_CE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(19[3:10])
    inout [15:0]SRAM_DATA;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(20[3:12])
    output [17:0]SRAM_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    input PIC_OE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(23[3:9])
    input PIC_WE_IN;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    input PIC_CS;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(25[3:9])
    input [18:0]PIC_ADDR_IN;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    inout [15:0]PIC_DATA_IN;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(27[3:14])
    output PIC_READY;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(28[3:12])
    output [7:0]LED;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    
    wire CLK_c /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    wire PIXEL_CLOCK /* synthesis SET_AS_NETWORK=PIXEL_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(43[8:19])
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(91[8:15])
    wire LOGIC_CLOCK_N_57 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    wire PIXEL_CLOCK_N_293 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(88[9:22])
    
    wire GND_net, VCC_net, Matrix_DATA_Out_c_11, Matrix_DATA_Out_c_10, 
        Matrix_DATA_Out_c_9, Matrix_DATA_Out_c_8, Matrix_DATA_Out_c_7, 
        Matrix_DATA_Out_c_6, Matrix_DATA_Out_c_5, Matrix_DATA_Out_c_4, 
        Matrix_DATA_Out_c_3, Matrix_DATA_Out_c_2, Matrix_DATA_Out_c_1, 
        Matrix_DATA_Out_c_0, Matrix_LINE_SEL_Out_c_2, Matrix_LINE_SEL_Out_c_1, 
        Matrix_LINE_SEL_Out_c_0, Matrix_CTRL_Out_c_2, Matrix_CTRL_Out_c_1, 
        Matrix_CTRL_Out_c_0, SRAM_OE_c, SRAM_WE_c, SRAM_ADDR_c_17, SRAM_ADDR_c_16, 
        SRAM_ADDR_c_15, SRAM_ADDR_c_14, SRAM_ADDR_c_13, SRAM_ADDR_c_12, 
        SRAM_ADDR_c_11, SRAM_ADDR_c_10, SRAM_ADDR_c_9, SRAM_ADDR_c_8, 
        SRAM_ADDR_c_7, SRAM_ADDR_c_6, SRAM_ADDR_c_5, SRAM_ADDR_c_4, 
        SRAM_ADDR_c_3, SRAM_ADDR_c_2, SRAM_ADDR_c_1, SRAM_ADDR_c_0, 
        PIC_OE_c, PIC_WE_IN_c, PIC_ADDR_IN_c_18, PIC_ADDR_IN_c_17, PIC_ADDR_IN_c_16, 
        PIC_ADDR_IN_c_15, PIC_ADDR_IN_c_14, PIC_ADDR_IN_c_13, PIC_ADDR_IN_c_12, 
        PIC_ADDR_IN_c_11, PIC_ADDR_IN_c_10, PIC_ADDR_IN_c_9, PIC_ADDR_IN_c_8, 
        PIC_ADDR_IN_c_7, PIC_ADDR_IN_c_6, PIC_ADDR_IN_c_5, PIC_ADDR_IN_c_4, 
        PIC_ADDR_IN_c_3, PIC_ADDR_IN_c_2, PIC_ADDR_IN_c_1, PIC_ADDR_IN_c_0, 
        PIC_READY_c;
    wire [15:0]BUS_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(48[8:16])
    wire [31:0]BUS_addr;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    wire [3:0]BUS_req;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(54[8:15])
    wire [3:0]BUS_currGrantID;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    wire [15:0]PIC_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(58[8:16])
    
    wire n15436, n4269;
    wire [15:0]MDM_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(73[8:16])
    
    wire n17458, n4575, n17457, n17456, BUS_DONE_OVERRIDE;
    wire [9:0]VRAM_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(88[8:17])
    wire [29:0]VRAM_DATA;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(89[8:17])
    wire [29:0]VRAM_DATA_OUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(90[8:21])
    
    wire VRAM_WE;
    wire [4:0]MATRIX_CURRROW;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(94[8:22])
    
    wire n4515, n17289, n17453, n4513, n17452, n4616, n4612, n4606, 
        n4602, n4618, n4617, BUS_currGrantID_3__N_55, n4260;
    wire [3:0]BUS_currGrantID_3__N_74;
    
    wire n40;
    wire [7:0]currPixel;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(65[9:18])
    wire [15:0]\PWMArray[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(79[9:17])
    
    wire n14080, SRAM_DATA_out_12, SRAM_DATA_out_11, n15469, SRAM_DATA_out_14, 
        SRAM_DATA_out_7;
    wire [15:0]currPWMCount;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(92[9:21])
    
    wire n4505, n4459;
    wire [15:0]currPWMCountMax;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(93[9:24])
    
    wire WRITE_DONE, n2877, n17272, n4611, n4581, n4601, n4595, 
        n4516, n4504, n4623, n14079, n14078, n14077, n14076, n14075, 
        n14074, n4460, n41, n6340;
    wire [7:0]state;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(87[9:14])
    
    wire n4397;
    wire [7:0]xOffset;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(96[9:16])
    wire [7:0]yOffset;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(97[9:16])
    
    wire n4498, n4306, n4307, n4508, n4304;
    wire [31:0]BUS_ADDR_INTERNAL;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(116[9:26])
    wire [15:0]otherData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(121[9:18])
    
    wire reset;
    wire [15:0]BUS_DATA_INTERNAL_adj_2580;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(128[9:26])
    wire [3:0]latchMode;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(145[9:18])
    
    wire SRAM_DATA_out_13, LOGIC_CLOCK_enable_52;
    wire [15:0]Sprite_readData2;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(174[9:25])
    
    wire n16341, n16340, n16338;
    wire [7:0]SpriteRead_yInSprite;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(185[9:29])
    wire [15:0]currSprite_size;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(194[9:24])
    
    wire n18264, n52;
    wire [8:0]RED_WRITE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(219[9:18])
    wire [8:0]GREEN_WRITE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(220[9:20])
    wire [8:0]BLUE_WRITE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(221[9:19])
    wire [8:0]ALPHA_WRITE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(222[9:20])
    
    wire SRAM_DATA_out_8, n4574, n16337, n16335, n16334, n16332, 
        n16331, n18263;
    wire [7:0]SpriteRead_yInSprite_7__N_597;
    wire [7:0]SpriteRead_yValid_N_1158;
    
    wire n51;
    wire [15:0]Sprite_readAddr_13__N_752;
    
    wire n4481, n4281, n59, n4560, state_7__N_345, n16329, n50, 
        n16328, n4503, n16326, n2801, n2802, n2803, n2804, n16325, 
        n4586, n4562, n4577, n4598, n8, n4596, LOGIC_CLOCK_N_57_enable_3, 
        n4376, n4559, n4374, n16321, n4387, n4373, n4372, n4371, 
        n4370, n16320, n4368, n4367, n4366, n4365, n4364, n4363, 
        n4394, n4558, n4557, n4476, n4597, n4613, n4615, n4593, 
        n4600, n4583, n4483, n4487, n4488, n4489, n4594, n4263, 
        n4259, n4264, n58, n4283, n4258, n1840, n4471, n4582, 
        n4604, n17287, n4614, n4592, n4591, n16316, n4, n16315, 
        n4496, n3296, n2642, n42, SRAM_DATA_out_9, n16313, n36, 
        n16312, n16310, n16309, n4295, n4294, n4293, n4292, n4291, 
        n4290, n4289, n4288, n4_adj_2523, n57, n49, n48, n4_adj_2524, 
        n4607, n16307, n16306, n16304, n16303, n16299, n4493, 
        n4494, n16298, n4509, n4390, n4389, n4388, n4452, n4453, 
        n4454, n4455, n4456, n4457, n4458, n4461, n4_adj_2525, 
        n16294, n16293, n16291, n16290, n4566, n4584, n4277, n16288, 
        n4470, n4517, n14, n16287, n16285, n4462, n18262, n4386, 
        n4385, n4384, n4393, n4621, n4619, n4490, n4265, n4620, 
        n4266, n4500, n16284, n16282, n16281, n16279, n16278, 
        n43, n16276, n16275, n4463, n4464, n4465, n4467, n17276, 
        n4480, n45, n46, n16271, n16270, n17434, n15771, n16266, 
        n4510, n16265, n4512, n4308, n4511, n4499, n16263, n4305, 
        n4247, n8_adj_2526, n4252, n4280, n4410, n4409, n4408, 
        n4407, n4406, n4405, n4404, n15539, n16262, n4299, n4298, 
        n4297, n4296, n4300, n4301, n16260, n16259, BUS_DONE_OUT_N_1051, 
        Sprite_pointers_N_1136, Sprite_pointers_N_1123, n4402, n4401, 
        n44, n16257, n16256, n16252, n4261, n16251, n4251, n4286, 
        n4362, n4466, n4272, n4608, n18261, n4_adj_2527, n4413, 
        n4412, n4250, n4248, n6, n16247, n4249, n4285, n16246, 
        n2504, n4475, n15770, n15768, n4603, n16244, n4479, n4268, 
        n4267, n4284, n4400, n4468, n4469, n16243, n16241, n4378, 
        n4377, n4256, n4605, n4570, n4565, n16240, n4403, n4568, 
        n16238, n4255, n4411, n4587, n17423, n16237, n4254, n16235, 
        n16234, n16232, n16231, n16223, n4474, n16222, n16221, 
        n47, n16220, n55, n16219, n56, n16218, n15767, n60, 
        n61, n33, n62;
    wire [31:0]lastAddress;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(29[8:19])
    wire [15:0]BUS_DATA_INTERNAL_adj_2601;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(30[8:25])
    
    wire BUS_DONE_INTERNAL, lastAddress_31__N_1328, lastAddress_31__N_1395, 
        lastAddress_31__N_1413, lastAddress_31__N_1333, lastAddress_31__N_1410, 
        lastAddress_31__N_1332, lastAddress_31__N_1407, lastAddress_31__N_1331, 
        lastAddress_31__N_1404, lastAddress_31__N_1330, lastAddress_31__N_1401, 
        lastAddress_31__N_1329, lastAddress_31__N_1398, lastAddress_31__N_1434, 
        lastAddress_31__N_1340, SRAM_WE_N_1254, n4563, n16217, n15765, 
        n16216, n6250, n4622, n4_adj_2532, n34, n2878, n63, n4572, 
        n15764, n4472, n4473, n15571, n4253, n64, n4478, n4477, 
        n4383, n4502, n4270, n4348, n4347, n15762, lastAddress_31__N_1310, 
        lastAddress_31__N_1327, lastAddress_31__N_1392, lastAddress_31__N_1326, 
        lastAddress_31__N_1389, lastAddress_31__N_1325, lastAddress_31__N_1386, 
        lastAddress_31__N_1324, lastAddress_31__N_1383, lastAddress_31__N_1323, 
        lastAddress_31__N_1380, lastAddress_31__N_1377, n15761, lastAddress_31__N_1431, 
        lastAddress_31__N_1339, lastAddress_31__N_1428, lastAddress_31__N_1338, 
        lastAddress_31__N_1425, lastAddress_31__N_1337, lastAddress_31__N_1422, 
        lastAddress_31__N_1336, lastAddress_31__N_1419, lastAddress_31__N_1335, 
        lastAddress_31__N_1416, lastAddress_31__N_1334, n16208, OUT_ENABLE, 
        BUS_DIRECTION_INTERNAL, n16207, n15759, n17275;
    wire [15:0]BUS_DATA_INTERNAL_adj_2609;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(39[8:25])
    
    wire n4352, n4353, n4354, n4391, n4356, n4357, n4358, n4359, 
        n4360, n4382;
    wire [31:0]BUS_ADDR_INTERNAL_adj_2610;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(40[8:25])
    
    wire WRITE_DONE_adj_2554, n4257;
    wire [15:0]writeData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(46[8:17])
    wire [7:0]state_adj_2613;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    
    wire n4350, n4514, n4375, n16206, n15758, n15756, n2880, n2879, 
        n4491, n16205, n16204, n4282, n4507, n4571, n16203, n4625, 
        n4396, n4369, n4588, n4495, n4501, n4482, n17411, n4361, 
        n16202, n4355, n16201, n39, n38, LOGIC_CLOCK_N_57_enable_7, 
        n4262, n17409, n4492, n4569, n4573, n4506, n4599, n10346, 
        n4287, n4278, n4243, n17408, n4567, n4271, n4242, n17407, 
        n4244, n4580, n4246, n4245, n4518, n4279, n4576, n4578, 
        n4579, n4585, n4590, n16497, n4610, n4564, n37, n4303, 
        n4273, n4302, n4609, n4392, n4395, n4351, n4497, n4399, 
        n4398, n16193, n16192, n4349, n35, n16191, n4561, n16190, 
        n16189, n16188, n16187, n16186, n63_adj_2556, n16178, n16177, 
        n15755, n16176, n15549, n15753, n16175, n16174, n63_adj_2557, 
        n15752, n15750, n15749, n15705, n16173, n16172, n16171, 
        LOGIC_CLOCK_N_57_enable_6, n15707, n16163, SRAM_DATA_out_10, 
        n16162, n16161, n14584, n16160, SRAM_DATA_out_15, SRAM_DATA_out_6, 
        SRAM_DATA_out_5, SRAM_DATA_out_4, SRAM_DATA_out_3, SRAM_DATA_out_2, 
        SRAM_DATA_out_1, SRAM_DATA_out_0, PIC_DATA_IN_out_15, PIC_DATA_IN_out_14, 
        PIC_DATA_IN_out_13, PIC_DATA_IN_out_12, PIC_DATA_IN_out_11, PIC_DATA_IN_out_10, 
        n16159, PIC_DATA_IN_out_9, PIC_DATA_IN_out_8, PIC_DATA_IN_out_7, 
        n16158, PIC_DATA_IN_out_6, PIC_DATA_IN_out_5, PIC_DATA_IN_out_4, 
        PIC_DATA_IN_out_3, n16157, PIC_DATA_IN_out_2, PIC_DATA_IN_out_1, 
        PIC_DATA_IN_out_0, n16156, n16456, n17394, n18278, n18277, 
        n4_adj_2558, n4_adj_2559, n18260, n16148, n16147, n16146, 
        n4_adj_2560, n16145, n16144, n16143, n15655, n16142, n16141, 
        n18280, n33_adj_2561, n16133, n16132, n16131, n16130, n4_adj_2562, 
        n16129, n15633, n17387, n16128, n16127, n9891, n16126, 
        n17385, n17384, n17383, n16122, n16121, n16115, n16114, 
        n17382, n17381, n16108, n16107, n18276, n18275, n16098, 
        n16097, n18274, n16085, n18273, n16084, n18272, n18271, 
        n18270, n18269, n13936, n5, n17380, n17379, n18268, n17378, 
        n17377, n18267, n18266, n18265, n17376, n17375, n17256, 
        n17374, n17373, BUS_ADDR_INTERNAL_18_derived_1, n17279, n17371, 
        n17368, n17366, n9950, n5_adj_2563, n17362, n17278, n17355, 
        n17274, n14_adj_2564, n9, n17344, n17343, n17342, n17340, 
        n17339, n15534, n17338, n18259, n17337, n17336, n17335, 
        n17334, n4_adj_2565, n17333, n9_adj_2566, n17332, n7, n17270, 
        n17331, n161, n17330, n17329, n160, n159, n13509, n17328, 
        n17327, n17326, n17325, n17323, n17322, n17321, n17320, 
        n5_adj_2567, n4_adj_2568, n17314, n17313, n17312, n17311, 
        n17310, n17309, n17308, n17307, n17305, n17304, n17302, 
        n17299, n17298;
    
    VHI i2 (.Z(VCC_net));
    BB SRAM_DATA_pad_11 (.I(BUS_data[11]), .T(SRAM_WE_c), .B(SRAM_DATA[11]), 
       .O(SRAM_DATA_out_11));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_5 (.I(BUS_data[5]), .T(SRAM_WE_c), .B(SRAM_DATA[5]), 
       .O(SRAM_DATA_out_5));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i3_4_lut (.A(PIC_data[0]), .B(n6), .C(\PWMArray[0] [9]), .D(n13509), 
         .Z(BUS_data[0])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i3_4_lut.init = 16'hfeee;
    LUT4 i2_4_lut (.A(BUS_DATA_INTERNAL_adj_2601[0]), .B(n17274), .C(n17330), 
         .D(BUS_DATA_INTERNAL_adj_2580[0]), .Z(n6)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i2_4_lut.init = 16'heca0;
    FD1P3DX BUS_currGrantID__i1 (.D(BUS_currGrantID_3__N_74[0]), .SP(LOGIC_CLOCK_N_57_enable_7), 
            .CK(LOGIC_CLOCK_N_57), .CD(BUS_currGrantID_3__N_55), .Q(BUS_currGrantID[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam BUS_currGrantID__i1.GSR = "DISABLED";
    LUT4 i12572_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4574), .D(n4558), 
         .Z(n16234)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12572_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12570_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4608), .D(n4592), 
         .Z(n16232)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12570_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12569_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4573), .D(n4557), 
         .Z(n16231)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12569_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12103_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4299), .D(n4283), 
         .Z(n15765)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12103_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12102_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4264), .D(n4248), 
         .Z(n15764)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12102_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12561_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4623), .D(n4607), 
         .Z(n16223)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12561_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12560_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4588), .D(n4572), 
         .Z(n16222)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12560_3_lut_4_lut.init = 16'hf4b0;
    SRAM RAM (.LOGIC_CLOCK(LOGIC_CLOCK), .lastAddress_31__N_1323(lastAddress_31__N_1323), 
         .n66({Open_0, n34, Open_1, Open_2, n37, n38, Open_3, 
         Open_4, Open_5, Open_6, Open_7, n44, Open_8, Open_9, 
         n47, n48, n49, n50, n51, n52, Open_10, Open_11, Open_12, 
         Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, 
         Open_20, Open_21}), .lastAddress_31__N_1386(lastAddress_31__N_1386), 
         .lastAddress_31__N_1324(lastAddress_31__N_1324), .lastAddress_31__N_1389(lastAddress_31__N_1389), 
         .lastAddress_31__N_1377(lastAddress_31__N_1377), .lastAddress_31__N_1310(lastAddress_31__N_1310), 
         .lastAddress_31__N_1325(lastAddress_31__N_1325), .lastAddress_31__N_1392(lastAddress_31__N_1392), 
         .lastAddress_31__N_1326(lastAddress_31__N_1326), .lastAddress_31__N_1395(lastAddress_31__N_1395), 
         .lastAddress_31__N_1327(lastAddress_31__N_1327), .lastAddress_31__N_1398(lastAddress_31__N_1398), 
         .BUS_DATA_INTERNAL({Open_22, Open_23, Open_24, Open_25, Open_26, 
         Open_27, Open_28, Open_29, Open_30, Open_31, Open_32, Open_33, 
         Open_34, Open_35, Open_36, BUS_DATA_INTERNAL_adj_2601[0]}), 
         .n17336(n17336), .SRAM_DATA_out_0(SRAM_DATA_out_0), .lastAddress_31__N_1328(lastAddress_31__N_1328), 
         .lastAddress_31__N_1401(lastAddress_31__N_1401), .lastAddress_31__N_1329(lastAddress_31__N_1329), 
         .lastAddress({Open_37, Open_38, Open_39, Open_40, Open_41, 
         Open_42, lastAddress[25], Open_43, Open_44, Open_45, Open_46, 
         Open_47, lastAddress[19:18], Open_48, Open_49, Open_50, Open_51, 
         Open_52, Open_53, Open_54, Open_55, Open_56, Open_57, Open_58, 
         lastAddress[6], Open_59, Open_60, Open_61, Open_62, Open_63, 
         lastAddress[0]}), .lastAddress_31__N_1410(lastAddress_31__N_1410), 
         .n56(n56), .SRAM_ADDR_c_0(SRAM_ADDR_c_0), .n17343(n17343), .lastAddress_31__N_1332(lastAddress_31__N_1332), 
         .n39(n39), .lastAddress_31__N_1339(lastAddress_31__N_1339), .lastAddress_31__N_1431(lastAddress_31__N_1431), 
         .n18280(n18280), .lastAddress_31__N_1380(lastAddress_31__N_1380), 
         .n46(n46), .lastAddress_31__N_1416(lastAddress_31__N_1416), .n58(n58), 
         .n45(n45), .lastAddress_31__N_1434(lastAddress_31__N_1434), .n64(n64), 
         .\BUS_ADDR_INTERNAL[18]_derived_1 (BUS_ADDR_INTERNAL_18_derived_1), 
         .lastAddress_31__N_1334(lastAddress_31__N_1334), .BUS_DONE_INTERNAL(BUS_DONE_INTERNAL), 
         .SRAM_WE_N_1254(SRAM_WE_N_1254), .\BUS_addr[10] (BUS_addr[10]), 
         .lastAddress_31__N_1404(lastAddress_31__N_1404), .\lastAddress[7] (lastAddress[7]), 
         .lastAddress_31__N_1413(lastAddress_31__N_1413), .n57(n57), .lastAddress_31__N_1419(lastAddress_31__N_1419), 
         .n59(n59), .n40(n40), .\lastAddress[5] (lastAddress[5]), .\lastAddress[24] (lastAddress[24]), 
         .SRAM_OE_c(SRAM_OE_c), .SRAM_WE_c(SRAM_WE_c), .lastAddress_31__N_1335(lastAddress_31__N_1335), 
         .n41(n41), .n18260(n18260), .n42(n42), .lastAddress_31__N_1422(lastAddress_31__N_1422), 
         .n60(n60), .n43(n43), .lastAddress_31__N_1340(lastAddress_31__N_1340), 
         .lastAddress_31__N_1336(lastAddress_31__N_1336), .n4(n4_adj_2532), 
         .\BUS_data[9] (BUS_data[9]), .\lastAddress[23] (lastAddress[23]), 
         .n4_adj_22(n4_adj_2523), .\BUS_data[10] (BUS_data[10]), .n4_adj_23(n4), 
         .\BUS_data[11] (BUS_data[11]), .n4_adj_24(n4_adj_2560), .\BUS_data[12] (BUS_data[12]), 
         .n4_adj_25(n4_adj_2559), .\BUS_data[13] (BUS_data[13]), .n4_adj_26(n4_adj_2558), 
         .\BUS_data[14] (BUS_data[14]), .lastAddress_31__N_1425(lastAddress_31__N_1425), 
         .n61(n61), .n4_adj_27(n4_adj_2527), .\BUS_data[15] (BUS_data[15]), 
         .\lastAddress[22] (lastAddress[22]), .n4_adj_28(n4_adj_2568), .\BUS_data[4] (BUS_data[4]), 
         .\lastAddress[4] (lastAddress[4]), .n4_adj_29(n4_adj_2524), .\BUS_data[5] (BUS_data[5]), 
         .n4_adj_30(n4_adj_2565), .\BUS_data[6] (BUS_data[6]), .lastAddress_31__N_1337(lastAddress_31__N_1337), 
         .n4_adj_31(n4_adj_2562), .\BUS_data[7] (BUS_data[7]), .lastAddress_31__N_1383(lastAddress_31__N_1383), 
         .lastAddress_31__N_1428(lastAddress_31__N_1428), .n62(n62), .\lastAddress[30] (lastAddress[30]), 
         .n33(n33), .n35(n35), .\lastAddress[21] (lastAddress[21]), .lastAddress_31__N_1338(lastAddress_31__N_1338), 
         .\BUS_DATA_INTERNAL[1] (BUS_DATA_INTERNAL_adj_2601[1]), .SRAM_DATA_out_1(SRAM_DATA_out_1), 
         .\BUS_DATA_INTERNAL[2] (BUS_DATA_INTERNAL_adj_2601[2]), .SRAM_DATA_out_2(SRAM_DATA_out_2), 
         .\BUS_DATA_INTERNAL[3] (BUS_DATA_INTERNAL_adj_2601[3]), .SRAM_DATA_out_3(SRAM_DATA_out_3), 
         .SRAM_DATA_out_4(SRAM_DATA_out_4), .SRAM_DATA_out_5(SRAM_DATA_out_5), 
         .SRAM_DATA_out_6(SRAM_DATA_out_6), .SRAM_DATA_out_7(SRAM_DATA_out_7), 
         .\BUS_DATA_INTERNAL[8] (BUS_DATA_INTERNAL_adj_2601[8]), .SRAM_DATA_out_8(SRAM_DATA_out_8), 
         .SRAM_DATA_out_9(SRAM_DATA_out_9), .SRAM_DATA_out_10(SRAM_DATA_out_10), 
         .SRAM_DATA_out_11(SRAM_DATA_out_11), .SRAM_DATA_out_12(SRAM_DATA_out_12), 
         .SRAM_DATA_out_13(SRAM_DATA_out_13), .SRAM_DATA_out_14(SRAM_DATA_out_14), 
         .SRAM_DATA_out_15(SRAM_DATA_out_15), .lastAddress_31__N_1333(lastAddress_31__N_1333), 
         .n36(n36), .\lastAddress[3] (lastAddress[3]), .\lastAddress[20] (lastAddress[20]), 
         .SRAM_ADDR_c_1(SRAM_ADDR_c_1), .n17342(n17342), .SRAM_ADDR_c_2(SRAM_ADDR_c_2), 
         .n17339(n17339), .SRAM_ADDR_c_3(SRAM_ADDR_c_3), .n17333(n17333), 
         .SRAM_ADDR_c_4(SRAM_ADDR_c_4), .n17332(n17332), .SRAM_ADDR_c_5(SRAM_ADDR_c_5), 
         .n17331(n17331), .SRAM_ADDR_c_6(SRAM_ADDR_c_6), .n17321(n17321), 
         .SRAM_ADDR_c_7(SRAM_ADDR_c_7), .n17334(n17334), .SRAM_ADDR_c_8(SRAM_ADDR_c_8), 
         .n17337(n17337), .SRAM_ADDR_c_9(SRAM_ADDR_c_9), .n17325(n17325), 
         .SRAM_ADDR_c_10(SRAM_ADDR_c_10), .SRAM_ADDR_c_11(SRAM_ADDR_c_11), 
         .\BUS_addr[11] (BUS_addr[11]), .SRAM_ADDR_c_12(SRAM_ADDR_c_12), 
         .n17335(n17335), .SRAM_ADDR_c_13(SRAM_ADDR_c_13), .n17338(n17338), 
         .SRAM_ADDR_c_14(SRAM_ADDR_c_14), .n17322(n17322), .SRAM_ADDR_c_15(SRAM_ADDR_c_15), 
         .n17320(n17320), .SRAM_ADDR_c_16(SRAM_ADDR_c_16), .n17323(n17323), 
         .SRAM_ADDR_c_17(SRAM_ADDR_c_17), .n17340(n17340), .lastAddress_31__N_1331(lastAddress_31__N_1331), 
         .lastAddress_31__N_1407(lastAddress_31__N_1407), .lastAddress_31__N_1330(lastAddress_31__N_1330), 
         .\lastAddress[2] (lastAddress[2]), .\lastAddress[31] (lastAddress[31]), 
         .n63(n63), .\lastAddress[17] (lastAddress[17]), .\lastAddress[29] (lastAddress[29]), 
         .\lastAddress[13] (lastAddress[13]), .\lastAddress[12] (lastAddress[12]), 
         .GND_net(GND_net), .\lastAddress[16] (lastAddress[16]), .\lastAddress[15] (lastAddress[15]), 
         .\lastAddress[14] (lastAddress[14]), .\lastAddress[28] (lastAddress[28]), 
         .\lastAddress[27] (lastAddress[27]), .\lastAddress[26] (lastAddress[26]), 
         .\lastAddress[1] (lastAddress[1]), .n55(n55), .\lastAddress[9] (lastAddress[9]), 
         .n17287(n17287), .n7(n7), .n9(n9_adj_2566), .n6250(n6250), 
         .\lastAddress[8] (lastAddress[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(199[7:23])
    BB SRAM_DATA_pad_6 (.I(BUS_data[6]), .T(SRAM_WE_c), .B(SRAM_DATA[6]), 
       .O(SRAM_DATA_out_6));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i12559_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4518), .D(n4502), 
         .Z(n16221)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12559_3_lut_4_lut.init = 16'hf4b0;
    MatrixDriver MD (.MATRIX_CURRROW({MATRIX_CURRROW}), .PIXEL_CLOCK(PIXEL_CLOCK), 
            .PIXEL_CLOCK_N_293(PIXEL_CLOCK_N_293), .WRITE_DONE(WRITE_DONE), 
            .LOGIC_CLOCK_N_57(LOGIC_CLOCK_N_57), .n18280(n18280), .currPWMCount({Open_64, 
            Open_65, Open_66, Open_67, Open_68, currPWMCount[10:7], 
            Open_69, Open_70, Open_71, Open_72, Open_73, Open_74, 
            currPWMCount[0]}), .LOGIC_CLOCK(LOGIC_CLOCK), .Matrix_CTRL_Out_c_1(Matrix_CTRL_Out_c_1), 
            .currPixel({currPixel}), .GND_net(GND_net), .Matrix_LINE_SEL_Out_c_1(Matrix_LINE_SEL_Out_c_1), 
            .n17305(n17305), .n17380(n17380), .n13509(n13509), .n15436(n15436), 
            .n17278(n17278), .n17373(n17373), .n18260(n18260), .\currPWMCountMax[1] (currPWMCountMax[1]), 
            .\currPWMCountMax[2] (currPWMCountMax[2]), .\currPWMCountMax[3] (currPWMCountMax[3]), 
            .\currPWMCountMax[4] (currPWMCountMax[4]), .\currPWMCountMax[5] (currPWMCountMax[5]), 
            .\currPWMCountMax[6] (currPWMCountMax[6]), .LOGIC_CLOCK_N_57_enable_6(LOGIC_CLOCK_N_57_enable_6), 
            .\BUS_data[3] (BUS_data[3]), .\currPWMCountMax[10] (currPWMCountMax[10]), 
            .\currPWMCountMax[12] (currPWMCountMax[12]), .\PWMArray[0][9] (\PWMArray[0] [9]), 
            .\currPWMCountMax[0] (currPWMCountMax[0]), .Matrix_LINE_SEL_Out_c_0(Matrix_LINE_SEL_Out_c_0), 
            .n17411(n17411), .n17458(n17458), .n16456(n16456), .n17368(n17368), 
            .\SpriteRead_yValid_N_1158[4] (SpriteRead_yValid_N_1158[4]), .n8(n8), 
            .n17371(n17371), .n17382(n17382), .n17374(n17374), .n17329(n17329), 
            .\currPWMCount[12] (currPWMCount[12]), .\currPWMCount[11] (currPWMCount[11]), 
            .\currPWMCount[6] (currPWMCount[6]), .\currPWMCount[5] (currPWMCount[5]), 
            .\currPWMCount[4] (currPWMCount[4]), .\currPWMCount[3] (currPWMCount[3]), 
            .\currPWMCount[2] (currPWMCount[2]), .\currPWMCount[1] (currPWMCount[1]), 
            .\BUS_data[2] (BUS_data[2]), .\BUS_data[0] (BUS_data[0]), .\BUS_data[1] (BUS_data[1]), 
            .\currPWMCountMax[11] (currPWMCountMax[11]), .\currPWMCountMax[9] (currPWMCountMax[9]), 
            .\currPWMCountMax[8] (currPWMCountMax[8]), .\currPWMCountMax[7] (currPWMCountMax[7]), 
            .n17326(n17326), .n17366(n17366), .n17407(n17407), .n17453(n17453), 
            .n17452(n17452), .\SpriteRead_yValid_N_1158[2] (SpriteRead_yValid_N_1158[2]), 
            .n15549(n15549), .n17289(n17289), .n17408(n17408), .\SpriteRead_yValid_N_1158[1] (SpriteRead_yValid_N_1158[1]), 
            .\SpriteRead_yValid_N_1158[0] (SpriteRead_yValid_N_1158[0]), .n4(n4_adj_2525), 
            .Matrix_CTRL_Out_c_2(Matrix_CTRL_Out_c_2), .n15705(n15705), 
            .n1840(n1840), .\BUS_currGrantID[0] (BUS_currGrantID[0]), .\BUS_currGrantID[1] (BUS_currGrantID[1]), 
            .\BUS_ADDR_INTERNAL[18] (BUS_ADDR_INTERNAL_adj_2610[18]), .lastAddress_31__N_1310(lastAddress_31__N_1310), 
            .\BUS_ADDR_INTERNAL[16] (BUS_ADDR_INTERNAL_adj_2610[16]), .n18277(n18277), 
            .\BUS_ADDR_INTERNAL[17] (BUS_ADDR_INTERNAL_adj_2610[17]), .n18264(n18264), 
            .\BUS_ADDR_INTERNAL[14] (BUS_ADDR_INTERNAL_adj_2610[14]), .n18262(n18262), 
            .\BUS_ADDR_INTERNAL[15] (BUS_ADDR_INTERNAL_adj_2610[15]), .n18271(n18271), 
            .n3296(n3296), .Matrix_DATA_Out_c_11(Matrix_DATA_Out_c_11), 
            .Matrix_DATA_Out_c_10(Matrix_DATA_Out_c_10), .Matrix_DATA_Out_c_9(Matrix_DATA_Out_c_9), 
            .Matrix_DATA_Out_c_8(Matrix_DATA_Out_c_8), .Matrix_DATA_Out_c_7(Matrix_DATA_Out_c_7), 
            .Matrix_DATA_Out_c_6(Matrix_DATA_Out_c_6), .Matrix_DATA_Out_c_5(Matrix_DATA_Out_c_5), 
            .\BUS_ADDR_INTERNAL[12] (BUS_ADDR_INTERNAL_adj_2610[12]), .n18272(n18272), 
            .\BUS_ADDR_INTERNAL[13] (BUS_ADDR_INTERNAL_adj_2610[13]), .n18266(n18266), 
            .Matrix_DATA_Out_c_4(Matrix_DATA_Out_c_4), .Matrix_DATA_Out_c_3(Matrix_DATA_Out_c_3), 
            .Matrix_DATA_Out_c_2(Matrix_DATA_Out_c_2), .\BUS_ADDR_INTERNAL[10] (BUS_ADDR_INTERNAL_adj_2610[10]), 
            .n18269(n18269), .\BUS_ADDR_INTERNAL[11] (BUS_ADDR_INTERNAL_adj_2610[11]), 
            .n18273(n18273), .\BUS_ADDR_INTERNAL[8] (BUS_ADDR_INTERNAL_adj_2610[8]), 
            .n18267(n18267), .\BUS_ADDR_INTERNAL[9] (BUS_ADDR_INTERNAL_adj_2610[9]), 
            .n18268(n18268), .\BUS_ADDR_INTERNAL[7] (BUS_ADDR_INTERNAL_adj_2610[7]), 
            .n18274(n18274), .Matrix_DATA_Out_c_1(Matrix_DATA_Out_c_1), 
            .Matrix_DATA_Out_c_0(Matrix_DATA_Out_c_0), .Matrix_LINE_SEL_Out_c_2(Matrix_LINE_SEL_Out_c_2), 
            .Matrix_CTRL_Out_c_0(Matrix_CTRL_Out_c_0), .\SpriteRead_yValid_N_1158[3] (SpriteRead_yValid_N_1158[3]), 
            .n17299(n17299), .\BUS_ADDR_INTERNAL[5] (BUS_ADDR_INTERNAL_adj_2610[5]), 
            .n18265(n18265), .\BUS_ADDR_INTERNAL[6] (BUS_ADDR_INTERNAL_adj_2610[6]), 
            .n18276(n18276), .\BUS_ADDR_INTERNAL[3] (BUS_ADDR_INTERNAL_adj_2610[3]), 
            .n17409(n17409), .\BUS_ADDR_INTERNAL[4] (BUS_ADDR_INTERNAL_adj_2610[4]), 
            .n18275(n18275), .\BUS_ADDR_INTERNAL[1] (BUS_ADDR_INTERNAL_adj_2610[1]), 
            .n17423(n17423), .\BUS_ADDR_INTERNAL[2] (BUS_ADDR_INTERNAL_adj_2610[2]), 
            .n18263(n18263), .\BUS_ADDR_INTERNAL[0] (BUS_ADDR_INTERNAL_adj_2610[0]), 
            .n18261(n18261), .\SpriteRead_yInSprite_7__N_597[0] (SpriteRead_yInSprite_7__N_597[0]), 
            .n17328(n17328), .n15539(n15539), .n17304(n17304), .n161(n161), 
            .n160(n160), .n159(n159), .n15633(n15633), .n17307(n17307), 
            .VRAM_DATA({VRAM_DATA}), .\VRAM_ADDR[8] (VRAM_ADDR[8]), .\VRAM_ADDR[7] (VRAM_ADDR[7]), 
            .\VRAM_ADDR[6] (VRAM_ADDR[6]), .\VRAM_ADDR[5] (VRAM_ADDR[5]), 
            .\VRAM_ADDR[4] (VRAM_ADDR[4]), .\VRAM_ADDR[3] (VRAM_ADDR[3]), 
            .\VRAM_ADDR[2] (VRAM_ADDR[2]), .\VRAM_ADDR[1] (VRAM_ADDR[1]), 
            .\VRAM_ADDR[0] (VRAM_ADDR[0]), .VRAM_WC(VRAM_WC), .VCC_net(VCC_net), 
            .VRAM_WE(VRAM_WE), .VRAM_DATA_OUT({VRAM_DATA_OUT}));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(142[6:30])
    LUT4 i12558_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4483), .D(n4467), 
         .Z(n16220)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12558_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12557_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4413), .D(n4397), 
         .Z(n16219)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12557_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12556_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4378), .D(n4362), 
         .Z(n16218)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12556_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i13116_4_lut (.A(n16497), .B(n17304), .C(n17373), .D(n17278), 
         .Z(LOGIC_CLOCK_N_57_enable_6)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i13116_4_lut.init = 16'h2000;
    LUT4 i12555_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4308), .D(n4292), 
         .Z(n16217)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12555_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12554_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4273), .D(n4257), 
         .Z(n16216)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12554_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6836_2_lut_rep_463 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL_adj_2610[1]), .Z(n18259)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam i6836_2_lut_rep_463.init = 16'h4040;
    LUT4 i12100_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4298), .D(n4282), 
         .Z(n15762)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12100_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12099_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4263), .D(n4247), 
         .Z(n15761)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12099_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12097_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4297), .D(n4281), 
         .Z(n15759)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12097_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12096_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4262), .D(n4246), 
         .Z(n15758)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12096_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_3_lut_rep_474 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(reset), .Z(n18270)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i1_2_lut_3_lut_rep_474.init = 16'h2020;
    LUT4 SRAM_WE_I_179_2_lut_rep_328_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(reset), .D(BUS_ADDR_INTERNAL_adj_2610[18]), 
         .Z(n17336)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam SRAM_WE_I_179_2_lut_rep_328_3_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i12094_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4296), .D(n4280), 
         .Z(n15756)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12094_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6648_2_lut_rep_335_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[0]), .D(BUS_ADDR_INTERNAL_adj_2610[0]), .Z(n17343)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6648_2_lut_rep_335_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i12093_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4261), .D(n4245), 
         .Z(n15755)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12093_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12091_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4295), .D(n4279), 
         .Z(n15753)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12091_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12090_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4260), .D(n4244), 
         .Z(n15752)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12090_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12546_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4622), .D(n4606), 
         .Z(n16208)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12546_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12545_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4587), .D(n4571), 
         .Z(n16207)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12545_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12544_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4517), .D(n4501), 
         .Z(n16206)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12544_3_lut_4_lut.init = 16'hf4b0;
    LUT4 SRAM_WE_N_1255_I_0_285_2_lut_3_lut_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(reset), .D(BUS_ADDR_INTERNAL_adj_2610[18]), 
         .Z(lastAddress_31__N_1377)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam SRAM_WE_N_1255_I_0_285_2_lut_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6420;
    LUT4 i12543_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4482), .D(n4466), 
         .Z(n16205)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12543_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12542_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4412), .D(n4396), 
         .Z(n16204)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12542_3_lut_4_lut.init = 16'hf4b0;
    LUT4 SRAM_WE_N_1255_I_0_286_2_lut_3_lut_4_lut_4_lut_3_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(reset), .Z(lastAddress_31__N_1380)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam SRAM_WE_N_1255_I_0_286_2_lut_3_lut_4_lut_4_lut_3_lut.init = 16'h2020;
    LUT4 i12541_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4377), .D(n4361), 
         .Z(n16203)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12541_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6799_2_lut_rep_466 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[14]), .Z(n18262)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6799_2_lut_rep_466.init = 16'h2020;
    LUT4 i12540_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4307), .D(n4291), 
         .Z(n16202)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12540_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12539_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4272), .D(n4256), 
         .Z(n16201)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12539_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12531_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4621), .D(n4605), 
         .Z(n16193)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12531_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12530_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4586), .D(n4570), 
         .Z(n16192)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12530_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12529_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4516), .D(n4500), 
         .Z(n16191)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12529_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6800_2_lut_rep_475 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[15]), .Z(n18271)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6800_2_lut_rep_475.init = 16'h2020;
    LUT4 i12528_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4481), .D(n4465), 
         .Z(n16190)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12528_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6900_2_lut_rep_312_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[15]), .D(BUS_ADDR_INTERNAL_adj_2610[15]), 
         .Z(n17320)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6900_2_lut_rep_312_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i12527_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4411), .D(n4395), 
         .Z(n16189)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12527_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6797_2_lut_rep_476 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[12]), .Z(n18272)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6797_2_lut_rep_476.init = 16'h2020;
    LUT4 i12526_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4376), .D(n4360), 
         .Z(n16188)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12526_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6899_2_lut_rep_314_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[14]), .D(BUS_ADDR_INTERNAL_adj_2610[14]), 
         .Z(n17322)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6899_2_lut_rep_314_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i12525_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4306), .D(n4290), 
         .Z(n16187)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12525_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12524_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4271), .D(n4255), 
         .Z(n16186)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12524_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12088_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4294), .D(n4278), 
         .Z(n15750)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12088_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6897_2_lut_rep_327_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[12]), .D(BUS_ADDR_INTERNAL_adj_2610[12]), 
         .Z(n17335)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6897_2_lut_rep_327_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i6796_2_lut_3_lut_rep_477 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[11]), .Z(n18273)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6796_2_lut_3_lut_rep_477.init = 16'h2020;
    LUT4 i12087_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4259), .D(n4243), 
         .Z(n15749)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12087_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6787_2_lut_rep_467 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[2]), .Z(n18263)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6787_2_lut_rep_467.init = 16'h2020;
    LUT4 i12516_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4620), .D(n4604), 
         .Z(n16178)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12516_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12515_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4585), .D(n4569), 
         .Z(n16177)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12515_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12514_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4515), .D(n4499), 
         .Z(n16176)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12514_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12513_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4480), .D(n4464), 
         .Z(n16175)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12513_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12512_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4410), .D(n4394), 
         .Z(n16174)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12512_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12511_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4375), .D(n4359), 
         .Z(n16173)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12511_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12510_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4305), .D(n4289), 
         .Z(n16172)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12510_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12509_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4270), .D(n4254), 
         .Z(n16171)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12509_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12501_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4619), .D(n4603), 
         .Z(n16163)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12501_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i2_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[11]), .D(BUS_ADDR_INTERNAL_adj_2610[11]), 
         .Z(BUS_addr[11])) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i2_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i12500_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4584), .D(n4568), 
         .Z(n16162)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12500_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12499_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4514), .D(n4498), 
         .Z(n16161)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12499_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12498_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4479), .D(n4463), 
         .Z(n16160)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12498_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12497_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4409), .D(n4393), 
         .Z(n16159)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12497_3_lut_4_lut.init = 16'hf4b0;
    FD1P3DX BUS_DONE_OVERRIDE_38 (.D(n18280), .SP(LOGIC_CLOCK_N_57_enable_3), 
            .CK(LOGIC_CLOCK_N_57), .CD(BUS_currGrantID_3__N_55), .Q(BUS_DONE_OVERRIDE)) /* synthesis lse_init_val=0 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam BUS_DONE_OVERRIDE_38.GSR = "DISABLED";
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i12496_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4374), .D(n4358), 
         .Z(n16158)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12496_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12495_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4304), .D(n4288), 
         .Z(n16157)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12495_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12494_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4269), .D(n4253), 
         .Z(n16156)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12494_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12486_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4618), .D(n4602), 
         .Z(n16148)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12486_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12485_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4583), .D(n4567), 
         .Z(n16147)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12485_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12484_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4513), .D(n4497), 
         .Z(n16146)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12484_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12483_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4478), .D(n4462), 
         .Z(n16145)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12483_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12482_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4408), .D(n4392), 
         .Z(n16144)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12482_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12481_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4373), .D(n4357), 
         .Z(n16143)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12481_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12480_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4303), .D(n4287), 
         .Z(n16142)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12480_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12479_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4268), .D(n4252), 
         .Z(n16141)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12479_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12471_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4617), .D(n4601), 
         .Z(n16133)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12471_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12470_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4582), .D(n4566), 
         .Z(n16132)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12470_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12469_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4512), .D(n4496), 
         .Z(n16131)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12469_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12468_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4477), .D(n4461), 
         .Z(n16130)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12468_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12467_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4407), .D(n4391), 
         .Z(n16129)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12467_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12466_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4372), .D(n4356), 
         .Z(n16128)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12466_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12465_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4302), .D(n4286), 
         .Z(n16127)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12465_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12464_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4267), .D(n4251), 
         .Z(n16126)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12464_3_lut_4_lut.init = 16'hf4b0;
    LUT4 lastAddress_i1_i15_3_lut_4_lut (.A(n17383), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[14]), .Z(n50)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i15_3_lut_4_lut.init = 16'hfb0b;
    LUT4 lastAddress_i1_i17_3_lut_4_lut (.A(n17362), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[16]), .Z(n48)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i17_3_lut_4_lut.init = 16'hfb0b;
    LUT4 lastAddress_i1_i10_3_lut_4_lut (.A(n17376), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[9]), .Z(n55)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i10_3_lut_4_lut.init = 16'hfb0b;
    BB SRAM_DATA_pad_12 (.I(BUS_data[12]), .T(SRAM_WE_c), .B(SRAM_DATA[12]), 
       .O(SRAM_DATA_out_12));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_7 (.I(BUS_data[7]), .T(SRAM_WE_c), .B(SRAM_DATA[7]), 
       .O(SRAM_DATA_out_7));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i6792_2_lut_rep_478 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[7]), .Z(n18274)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6792_2_lut_rep_478.init = 16'h2020;
    LUT4 lastAddress_i1_i6_3_lut_4_lut (.A(n17380), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[5]), .Z(n59)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i6_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i3_4_lut_adj_673 (.A(BUS_DONE_INTERNAL), .B(BUS_DONE_OVERRIDE), 
         .C(BUS_ADDR_INTERNAL_18_derived_1), .D(WRITE_DONE), .Z(n8_adj_2526)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:83])
    defparam i3_4_lut_adj_673.init = 16'hffce;
    BB SRAM_DATA_pad_8 (.I(BUS_data[8]), .T(SRAM_WE_c), .B(SRAM_DATA[8]), 
       .O(SRAM_DATA_out_8));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_13 (.I(BUS_data[13]), .T(SRAM_WE_c), .B(SRAM_DATA[13]), 
       .O(SRAM_DATA_out_13));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_14 (.I(BUS_data[14]), .T(SRAM_WE_c), .B(SRAM_DATA[14]), 
       .O(SRAM_DATA_out_14));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_10 (.I(BUS_data[10]), .T(SRAM_WE_c), .B(SRAM_DATA[10]), 
       .O(SRAM_DATA_out_10));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_9 (.I(BUS_data[9]), .T(SRAM_WE_c), .B(SRAM_DATA[9]), 
       .O(SRAM_DATA_out_9));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i6892_2_lut_rep_326_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[7]), .D(BUS_ADDR_INTERNAL_adj_2610[7]), .Z(n17334)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6892_2_lut_rep_326_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i6789_2_lut_rep_479 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[4]), .Z(n18275)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6789_2_lut_rep_479.init = 16'h2020;
    LUT4 lastAddress_i1_i5_3_lut_4_lut (.A(n17375), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[4]), .Z(n60)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i5_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_2_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[4]), .D(BUS_ADDR_INTERNAL_adj_2610[4]), .Z(n15436)) /* synthesis lut_function=(A (B+!(C))+!A !((D)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i1_2_lut_4_lut_4_lut_4_lut.init = 16'h8ace;
    LUT4 i6886_2_lut_rep_334_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(BUS_ADDR_INTERNAL_adj_2610[1]), .D(BUS_ADDR_INTERNAL[1]), 
         .Z(n17342)) /* synthesis lut_function=(!(A (B+!(D))+!A !((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam i6886_2_lut_rep_334_3_lut_4_lut_4_lut_4_lut.init = 16'h7351;
    LUT4 i6889_2_lut_rep_324_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[4]), .D(BUS_ADDR_INTERNAL_adj_2610[4]), .Z(n17332)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6889_2_lut_rep_324_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 lastAddress_i1_i4_3_lut_4_lut (.A(n17371), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[3]), .Z(n61)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i4_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i6791_2_lut_rep_480 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[6]), .Z(n18276)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6791_2_lut_rep_480.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n17373), .B(n17458), .C(Sprite_pointers_N_1123), 
         .D(n17374), .Z(n4625)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i6891_2_lut_rep_313_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[6]), .D(BUS_ADDR_INTERNAL_adj_2610[6]), .Z(n17321)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6891_2_lut_rep_313_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i6801_2_lut_rep_481 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[16]), .Z(n18277)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6801_2_lut_rep_481.init = 16'h2020;
    LUT4 i6887_2_lut_rep_331_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[2]), .D(BUS_ADDR_INTERNAL_adj_2610[2]), .Z(n17339)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6887_2_lut_rep_331_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_674 (.A(n17373), .B(n17458), .C(Sprite_pointers_N_1123), 
         .D(n17374), .Z(n4591)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_674.init = 16'h4000;
    LUT4 i6901_2_lut_rep_315_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[16]), .D(BUS_ADDR_INTERNAL_adj_2610[16]), 
         .Z(n17323)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6901_2_lut_rep_315_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 lastAddress_i1_i8_3_lut_4_lut (.A(n17373), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[7]), .Z(n57)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i8_3_lut_4_lut.init = 16'hfb0b;
    LUT4 PIC_dir_I_0_3_lut_rep_464 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_DIRECTION_INTERNAL), .Z(n18260)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam PIC_dir_I_0_3_lut_rep_464.init = 16'h6262;
    LUT4 i6802_2_lut_rep_468 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[17]), .Z(n18264)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6802_2_lut_rep_468.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n17373), .B(n17458), .C(Sprite_pointers_N_1123), 
         .D(n17374), .Z(n4590)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_332_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[17]), .D(BUS_ADDR_INTERNAL_adj_2610[17]), 
         .Z(n17340)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i1_2_lut_rep_332_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i6790_2_lut_rep_469 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[5]), .Z(n18265)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6790_2_lut_rep_469.init = 16'h2020;
    LUT4 lastAddress_i1_i13_3_lut_4_lut (.A(n17377), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[12]), .Z(n52)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i13_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_4_lut_4_lut_4_lut_rep_482 (.A(BUS_DIRECTION_INTERNAL), .B(BUS_currGrantID[0]), 
         .C(BUS_currGrantID[1]), .Z(n18278)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(107[13:31])
    defparam i1_4_lut_4_lut_4_lut_rep_482.init = 16'h1010;
    LUT4 i6890_2_lut_rep_323_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[5]), .D(BUS_ADDR_INTERNAL_adj_2610[5]), .Z(n17331)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6890_2_lut_rep_323_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i6968_2_lut_4_lut (.A(BUS_DIRECTION_INTERNAL), .B(BUS_currGrantID[0]), 
         .C(BUS_currGrantID[1]), .D(writeData[8]), .Z(PIC_data[8])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(107[13:31])
    defparam i6968_2_lut_4_lut.init = 16'h1000;
    LUT4 BUS_VALID_I_0_2_lut_rep_322_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(BUS_DIRECTION_INTERNAL), .D(BUS_ADDR_INTERNAL_adj_2610[18]), 
         .Z(n17330)) /* synthesis lut_function=(!(A (B)+!A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam BUS_VALID_I_0_2_lut_rep_322_3_lut_4_lut_4_lut_4_lut.init = 16'h2262;
    LUT4 i6798_2_lut_rep_470 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[13]), .Z(n18266)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6798_2_lut_rep_470.init = 16'h2020;
    LUT4 i6898_2_lut_rep_330_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[13]), .D(BUS_ADDR_INTERNAL_adj_2610[13]), 
         .Z(n17338)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6898_2_lut_rep_330_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i6582_2_lut_rep_465 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[0]), .Z(n18261)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6582_2_lut_rep_465.init = 16'h2020;
    LUT4 i6793_2_lut_rep_471 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[8]), .Z(n18267)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6793_2_lut_rep_471.init = 16'h2020;
    LUT4 i6893_2_lut_rep_329_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[8]), .D(BUS_ADDR_INTERNAL_adj_2610[8]), .Z(n17337)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6893_2_lut_rep_329_4_lut_4_lut_4_lut.init = 16'h7531;
    BB SRAM_DATA_pad_4 (.I(BUS_data[4]), .T(SRAM_WE_c), .B(SRAM_DATA[4]), 
       .O(SRAM_DATA_out_4));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i6794_2_lut_rep_472 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[9]), .Z(n18268)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6794_2_lut_rep_472.init = 16'h2020;
    BB SRAM_DATA_pad_15 (.I(BUS_data[15]), .T(SRAM_WE_c), .B(SRAM_DATA[15]), 
       .O(SRAM_DATA_out_15));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_3 (.I(BUS_data[3]), .T(SRAM_WE_c), .B(SRAM_DATA[3]), 
       .O(SRAM_DATA_out_3));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_2 (.I(BUS_data[2]), .T(SRAM_WE_c), .B(SRAM_DATA[2]), 
       .O(SRAM_DATA_out_2));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_1 (.I(BUS_data[1]), .T(SRAM_WE_c), .B(SRAM_DATA[1]), 
       .O(SRAM_DATA_out_1));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_0 (.I(BUS_data[0]), .T(SRAM_WE_c), .B(SRAM_DATA[0]), 
       .O(SRAM_DATA_out_0));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB PIC_DATA_IN_pad_15 (.I(BUS_data[15]), .T(PIC_OE_c), .B(PIC_DATA_IN[15]), 
       .O(PIC_DATA_IN_out_15));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_14 (.I(BUS_data[14]), .T(PIC_OE_c), .B(PIC_DATA_IN[14]), 
       .O(PIC_DATA_IN_out_14));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_13 (.I(BUS_data[13]), .T(PIC_OE_c), .B(PIC_DATA_IN[13]), 
       .O(PIC_DATA_IN_out_13));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_12 (.I(BUS_data[12]), .T(PIC_OE_c), .B(PIC_DATA_IN[12]), 
       .O(PIC_DATA_IN_out_12));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_11 (.I(BUS_data[11]), .T(PIC_OE_c), .B(PIC_DATA_IN[11]), 
       .O(PIC_DATA_IN_out_11));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_10 (.I(BUS_data[10]), .T(PIC_OE_c), .B(PIC_DATA_IN[10]), 
       .O(PIC_DATA_IN_out_10));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_9 (.I(BUS_data[9]), .T(PIC_OE_c), .B(PIC_DATA_IN[9]), 
       .O(PIC_DATA_IN_out_9));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_8 (.I(BUS_data[8]), .T(PIC_OE_c), .B(PIC_DATA_IN[8]), 
       .O(PIC_DATA_IN_out_8));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_7 (.I(BUS_data[7]), .T(PIC_OE_c), .B(PIC_DATA_IN[7]), 
       .O(PIC_DATA_IN_out_7));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_6 (.I(BUS_data[6]), .T(PIC_OE_c), .B(PIC_DATA_IN[6]), 
       .O(PIC_DATA_IN_out_6));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_5 (.I(BUS_data[5]), .T(PIC_OE_c), .B(PIC_DATA_IN[5]), 
       .O(PIC_DATA_IN_out_5));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_4 (.I(BUS_data[4]), .T(PIC_OE_c), .B(PIC_DATA_IN[4]), 
       .O(PIC_DATA_IN_out_4));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_3 (.I(BUS_data[3]), .T(PIC_OE_c), .B(PIC_DATA_IN[3]), 
       .O(PIC_DATA_IN_out_3));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_2 (.I(BUS_data[2]), .T(PIC_OE_c), .B(PIC_DATA_IN[2]), 
       .O(PIC_DATA_IN_out_2));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_1 (.I(BUS_data[1]), .T(PIC_OE_c), .B(PIC_DATA_IN[1]), 
       .O(PIC_DATA_IN_out_1));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_0 (.I(BUS_data[0]), .T(PIC_OE_c), .B(PIC_DATA_IN[0]), 
       .O(PIC_DATA_IN_out_0));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    OB UART_TX_pad (.I(GND_net), .O(UART_TX));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(11[3:10])
    OB Matrix_DATA_Out_pad_11 (.I(Matrix_DATA_Out_c_11), .O(Matrix_DATA_Out[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_10 (.I(Matrix_DATA_Out_c_10), .O(Matrix_DATA_Out[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_9 (.I(Matrix_DATA_Out_c_9), .O(Matrix_DATA_Out[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_8 (.I(Matrix_DATA_Out_c_8), .O(Matrix_DATA_Out[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_7 (.I(Matrix_DATA_Out_c_7), .O(Matrix_DATA_Out[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_6 (.I(Matrix_DATA_Out_c_6), .O(Matrix_DATA_Out[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_5 (.I(Matrix_DATA_Out_c_5), .O(Matrix_DATA_Out[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_4 (.I(Matrix_DATA_Out_c_4), .O(Matrix_DATA_Out[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_3 (.I(Matrix_DATA_Out_c_3), .O(Matrix_DATA_Out[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_2 (.I(Matrix_DATA_Out_c_2), .O(Matrix_DATA_Out[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_1 (.I(Matrix_DATA_Out_c_1), .O(Matrix_DATA_Out[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_0 (.I(Matrix_DATA_Out_c_0), .O(Matrix_DATA_Out[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_LINE_SEL_Out_pad_3 (.I(GND_net), .O(Matrix_LINE_SEL_Out[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_LINE_SEL_Out_pad_2 (.I(Matrix_LINE_SEL_Out_c_2), .O(Matrix_LINE_SEL_Out[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_LINE_SEL_Out_pad_1 (.I(Matrix_LINE_SEL_Out_c_1), .O(Matrix_LINE_SEL_Out[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_LINE_SEL_Out_pad_0 (.I(Matrix_LINE_SEL_Out_c_0), .O(Matrix_LINE_SEL_Out[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_CTRL_Out_pad_2 (.I(Matrix_CTRL_Out_c_2), .O(Matrix_CTRL_Out[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    OB Matrix_CTRL_Out_pad_1 (.I(Matrix_CTRL_Out_c_1), .O(Matrix_CTRL_Out[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    OB Matrix_CTRL_Out_pad_0 (.I(Matrix_CTRL_Out_c_0), .O(Matrix_CTRL_Out[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    OB SRAM_OE_pad (.I(SRAM_OE_c), .O(SRAM_OE));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(17[3:10])
    OB SRAM_WE_pad (.I(SRAM_WE_c), .O(SRAM_WE));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(18[3:10])
    OB SRAM_CE_pad (.I(GND_net), .O(SRAM_CE));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(19[3:10])
    OB SRAM_ADDR_pad_17 (.I(SRAM_ADDR_c_17), .O(SRAM_ADDR[17]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_16 (.I(SRAM_ADDR_c_16), .O(SRAM_ADDR[16]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_15 (.I(SRAM_ADDR_c_15), .O(SRAM_ADDR[15]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_14 (.I(SRAM_ADDR_c_14), .O(SRAM_ADDR[14]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_13 (.I(SRAM_ADDR_c_13), .O(SRAM_ADDR[13]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_12 (.I(SRAM_ADDR_c_12), .O(SRAM_ADDR[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_11 (.I(SRAM_ADDR_c_11), .O(SRAM_ADDR[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_10 (.I(SRAM_ADDR_c_10), .O(SRAM_ADDR[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_9 (.I(SRAM_ADDR_c_9), .O(SRAM_ADDR[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_8 (.I(SRAM_ADDR_c_8), .O(SRAM_ADDR[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_7 (.I(SRAM_ADDR_c_7), .O(SRAM_ADDR[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_6 (.I(SRAM_ADDR_c_6), .O(SRAM_ADDR[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_5 (.I(SRAM_ADDR_c_5), .O(SRAM_ADDR[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_4 (.I(SRAM_ADDR_c_4), .O(SRAM_ADDR[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_3 (.I(SRAM_ADDR_c_3), .O(SRAM_ADDR[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_2 (.I(SRAM_ADDR_c_2), .O(SRAM_ADDR[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_1 (.I(SRAM_ADDR_c_1), .O(SRAM_ADDR[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_0 (.I(SRAM_ADDR_c_0), .O(SRAM_ADDR[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB PIC_READY_pad (.I(PIC_READY_c), .O(PIC_READY));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(28[3:12])
    OB LED_pad_7 (.I(GND_net), .O(LED[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_6 (.I(GND_net), .O(LED[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_5 (.I(GND_net), .O(LED[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_4 (.I(GND_net), .O(LED[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_3 (.I(GND_net), .O(LED[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_2 (.I(GND_net), .O(LED[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_1 (.I(GND_net), .O(LED[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_0 (.I(GND_net), .O(LED[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    IB CLK_pad (.I(CLK), .O(CLK_c));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    IB PIC_OE_pad (.I(PIC_OE), .O(PIC_OE_c));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(23[3:9])
    IB PIC_WE_IN_pad (.I(PIC_WE_IN), .O(PIC_WE_IN_c));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    IB PIC_ADDR_IN_pad_18 (.I(PIC_ADDR_IN[18]), .O(PIC_ADDR_IN_c_18));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_17 (.I(PIC_ADDR_IN[17]), .O(PIC_ADDR_IN_c_17));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_16 (.I(PIC_ADDR_IN[16]), .O(PIC_ADDR_IN_c_16));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_15 (.I(PIC_ADDR_IN[15]), .O(PIC_ADDR_IN_c_15));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_14 (.I(PIC_ADDR_IN[14]), .O(PIC_ADDR_IN_c_14));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_13 (.I(PIC_ADDR_IN[13]), .O(PIC_ADDR_IN_c_13));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_12 (.I(PIC_ADDR_IN[12]), .O(PIC_ADDR_IN_c_12));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_11 (.I(PIC_ADDR_IN[11]), .O(PIC_ADDR_IN_c_11));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_10 (.I(PIC_ADDR_IN[10]), .O(PIC_ADDR_IN_c_10));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_9 (.I(PIC_ADDR_IN[9]), .O(PIC_ADDR_IN_c_9));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_8 (.I(PIC_ADDR_IN[8]), .O(PIC_ADDR_IN_c_8));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_7 (.I(PIC_ADDR_IN[7]), .O(PIC_ADDR_IN_c_7));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_6 (.I(PIC_ADDR_IN[6]), .O(PIC_ADDR_IN_c_6));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_5 (.I(PIC_ADDR_IN[5]), .O(PIC_ADDR_IN_c_5));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_4 (.I(PIC_ADDR_IN[4]), .O(PIC_ADDR_IN_c_4));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_3 (.I(PIC_ADDR_IN[3]), .O(PIC_ADDR_IN_c_3));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_2 (.I(PIC_ADDR_IN[2]), .O(PIC_ADDR_IN_c_2));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_1 (.I(PIC_ADDR_IN[1]), .O(PIC_ADDR_IN_c_1));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_0 (.I(PIC_ADDR_IN[0]), .O(PIC_ADDR_IN_c_0));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    LUT4 i13053_2_lut_rep_448 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .Z(n17456)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i13053_2_lut_rep_448.init = 16'h2222;
    FD1P3DX BUS_currGrantID__i2 (.D(BUS_currGrantID_3__N_74[1]), .SP(LOGIC_CLOCK_N_57_enable_7), 
            .CK(LOGIC_CLOCK_N_57), .CD(BUS_currGrantID_3__N_55), .Q(BUS_currGrantID[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam BUS_currGrantID__i2.GSR = "DISABLED";
    LUT4 i6786_2_lut_rep_415_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[1]), .Z(n17423)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6786_2_lut_rep_415_3_lut.init = 16'h2020;
    LUT4 i6788_2_lut_rep_401_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[3]), .Z(n17409)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6788_2_lut_rep_401_3_lut.init = 16'h2020;
    LUT4 n10147_bdd_2_lut_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(state[1]), .Z(n17256)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam n10147_bdd_2_lut_3_lut.init = 16'h0d0d;
    LUT4 lastAddress_i1_i9_3_lut_4_lut (.A(n17378), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[8]), .Z(n56)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i9_3_lut_4_lut.init = 16'hfb0b;
    LUT4 lastAddress_i1_i14_3_lut_4_lut (.A(n17379), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[13]), .Z(n51)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i14_3_lut_4_lut.init = 16'hfb0b;
    GSR GSR_INST (.GSR(state_7__N_345));
    LUT4 lastAddress_i1_i3_3_lut_4_lut (.A(n17382), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[2]), .Z(n62)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i3_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_2_lut_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(state[3]), .Z(n33_adj_2561)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i1_2_lut_3_lut.init = 16'hd0d0;
    LUT4 lastAddress_i1_i18_3_lut_4_lut (.A(n17458), .B(n17381), .C(SRAM_WE_N_1254), 
         .D(lastAddress[17]), .Z(n47)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam lastAddress_i1_i18_3_lut_4_lut.init = 16'hfd0d;
    LUT4 i10609_4_lut_4_lut (.A(n17458), .B(n17381), .C(n13936), .D(n17411), 
         .Z(BUS_DONE_OUT_N_1051)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i10609_4_lut_4_lut.init = 16'hfd55;
    LUT4 i6561_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(state[1]), .D(state[0]), .Z(n9891)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (C+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6561_3_lut_4_lut.init = 16'hffd0;
    LUT4 lastAddress_i1_i2_3_lut_4_lut (.A(n17384), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[1]), .Z(n63)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i2_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_783_i4_3_lut_4_lut (.A(n17384), .B(n17458), .C(latchMode[3]), 
         .D(n2801), .Z(n2877)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_783_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_783_i3_3_lut_4_lut (.A(n17384), .B(n17458), .C(latchMode[2]), 
         .D(n2802), .Z(n2878)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_783_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_783_i2_3_lut_4_lut (.A(n17384), .B(n17458), .C(latchMode[1]), 
         .D(n2803), .Z(n2879)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_783_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 equal_1134_i3_2_lut_rep_449 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .Z(n17457)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam equal_1134_i3_2_lut_rep_449.init = 16'hbbbb;
    LUT4 mux_783_i1_3_lut_4_lut (.A(n17384), .B(n17458), .C(latchMode[0]), 
         .D(n2804), .Z(n2880)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_783_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_GRANT_I_0_317_2_lut_rep_262_2_lut_3_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(n17275), .Z(n17270)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam BUS_GRANT_I_0_317_2_lut_rep_262_2_lut_3_lut.init = 16'h0404;
    LUT4 i1891_4_lut (.A(currPixel[7]), .B(currPixel[0]), .C(n15707), 
         .D(n17289), .Z(n1840)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(65[9:18])
    defparam i1891_4_lut.init = 16'h5f5d;
    LUT4 i12046_2_lut (.A(currPixel[1]), .B(n15705), .Z(n15707)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12046_2_lut.init = 16'heeee;
    LUT4 i12044_4_lut (.A(currPixel[3]), .B(currPixel[6]), .C(currPixel[5]), 
         .D(n15633), .Z(n15705)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12044_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n17385), .B(n17458), .C(n6340), 
         .D(n17384), .Z(n63_adj_2557)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i2_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'hfbff;
    LUT4 mux_767_i4_3_lut_4_lut (.A(n17385), .B(n17458), .C(yOffset[3]), 
         .D(xOffset[3]), .Z(n2801)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_767_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6853_2_lut_rep_403_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL_adj_2610[18]), .Z(n17411)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam i6853_2_lut_rep_403_3_lut.init = 16'h4040;
    LUT4 i11922_2_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(state_adj_2613[4]), .D(n17275), .Z(n14)) /* synthesis lut_function=(!(A (C)+!A (B (C (D))+!B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam i11922_2_lut_3_lut_3_lut_4_lut.init = 16'h0f4f;
    LUT4 i12422_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[5]), 
         .D(RED_WRITE[5]), .Z(n16084)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12422_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12423_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[5]), 
         .D(BLUE_WRITE[5]), .Z(n16085)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12423_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12435_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[1]), 
         .D(RED_WRITE[1]), .Z(n16097)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12435_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12436_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[1]), 
         .D(BLUE_WRITE[1]), .Z(n16098)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12436_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12445_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[6]), 
         .D(RED_WRITE[6]), .Z(n16107)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12445_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12446_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[6]), 
         .D(BLUE_WRITE[6]), .Z(n16108)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12446_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_DIRECTION_IN_I_0_1_lut_rep_379_3_lut_4_lut_3_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(BUS_DIRECTION_INTERNAL), .Z(n17387)) /* synthesis lut_function=(A (B)+!A !(B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam BUS_DIRECTION_IN_I_0_1_lut_rep_379_3_lut_4_lut_3_lut.init = 16'h9d9d;
    LUT4 i6616_2_lut_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_DIRECTION_INTERNAL), .Z(n9950)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(100[26:48])
    defparam i6616_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(n17385), .B(n17458), .C(n6340), 
         .D(n17384), .Z(n63_adj_2556)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i12608_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[2]), 
         .D(RED_WRITE[2]), .Z(n16270)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12608_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12609_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[2]), 
         .D(BLUE_WRITE[2]), .Z(n16271)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12609_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12636_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[3]), 
         .D(RED_WRITE[3]), .Z(n16298)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12636_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12637_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[3]), 
         .D(BLUE_WRITE[3]), .Z(n16299)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12637_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_450 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .Z(n17458)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i1_2_lut_rep_450.init = 16'heeee;
    LUT4 lastAddress_i1_i31_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[30]), .Z(n34)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i31_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i26_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[25]), .Z(n39)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i26_3_lut_4_lut.init = 16'hf101;
    LUT4 i13080_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_currGrantID_3__N_74[0]), .D(BUS_req[2]), .Z(LOGIC_CLOCK_N_57_enable_7)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i13080_3_lut_4_lut.init = 16'h1110;
    LUT4 i12658_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[4]), 
         .D(RED_WRITE[4]), .Z(n16320)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12658_3_lut_4_lut.init = 16'hf4b0;
    LUT4 lastAddress_i1_i21_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[20]), .Z(n44)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i21_3_lut_4_lut.init = 16'hf101;
    LUT4 i12659_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[4]), 
         .D(BLUE_WRITE[4]), .Z(n16321)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12659_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12460_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[8]), 
         .D(BLUE_WRITE[8]), .Z(n16122)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12460_3_lut_4_lut.init = 16'hf4b0;
    LUT4 lastAddress_i1_i27_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[26]), .Z(n38)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i27_3_lut_4_lut.init = 16'hf101;
    LUT4 i12589_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[0]), 
         .D(RED_WRITE[0]), .Z(n16251)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12589_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12590_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[0]), 
         .D(BLUE_WRITE[0]), .Z(n16252)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12590_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12452_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[7]), 
         .D(RED_WRITE[7]), .Z(n16114)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12452_3_lut_4_lut.init = 16'hf4b0;
    LUT4 lastAddress_i1_i28_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[27]), .Z(n37)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i28_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i20_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[19]), .Z(n45)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i20_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i25_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(SRAM_WE_N_1254), .D(lastAddress[24]), .Z(n40)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i25_3_lut_4_lut.init = 16'hf101;
    LUT4 i6742_3_lut_rep_319_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(n17373), .D(n17374), .Z(n17327)) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i6742_3_lut_rep_319_4_lut.init = 16'hf111;
    LUT4 i12453_3_lut_4_lut (.A(n17385), .B(n17458), .C(ALPHA_WRITE[7]), 
         .D(BLUE_WRITE[7]), .Z(n16115)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12453_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12459_3_lut_4_lut (.A(n17385), .B(n17458), .C(GREEN_WRITE[8]), 
         .D(RED_WRITE[8]), .Z(n16121)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12459_3_lut_4_lut.init = 16'hf4b0;
    LUT4 lastAddress_i1_i1_3_lut_4_lut (.A(n17385), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[0]), .Z(n64)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i1_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_767_i2_3_lut_4_lut (.A(n17385), .B(n17458), .C(yOffset[1]), 
         .D(xOffset[1]), .Z(n2803)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_767_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_767_i3_3_lut_4_lut (.A(n17385), .B(n17458), .C(yOffset[2]), 
         .D(xOffset[2]), .Z(n2802)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_767_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_767_i1_3_lut_4_lut (.A(n17385), .B(n17458), .C(yOffset[0]), 
         .D(xOffset[0]), .Z(n2804)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam mux_767_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i3212_3_lut_rep_306_4_lut (.A(n17362), .B(n17381), .C(n17411), 
         .D(n17458), .Z(n17314)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i3212_3_lut_rep_306_4_lut.init = 16'he0ff;
    LUT4 i1_2_lut_rep_301_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(n17374), .D(n17373), .Z(n17309)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i1_2_lut_rep_301_3_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i6772_2_lut_rep_305_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(n17374), .D(n17373), .Z(n17313)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i6772_2_lut_rep_305_3_lut_4_lut.init = 16'hfff1;
    CCU2D sub_991_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14080), .S0(n3296));
    defparam sub_991_add_2_cout.INIT0 = 16'h0000;
    defparam sub_991_add_2_cout.INIT1 = 16'h0000;
    defparam sub_991_add_2_cout.INJECT1_0 = "NO";
    defparam sub_991_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_991_add_2_13 (.A0(currPWMCount[11]), .B0(currPWMCountMax[11]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[12]), .B1(currPWMCountMax[12]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14079), .COUT(n14080));
    defparam sub_991_add_2_13.INIT0 = 16'h5999;
    defparam sub_991_add_2_13.INIT1 = 16'h5999;
    defparam sub_991_add_2_13.INJECT1_0 = "NO";
    defparam sub_991_add_2_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_300_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(n17374), .D(n17373), .Z(n17308)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i1_2_lut_rep_300_3_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i11996_2_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_addr[11]), .D(n17382), .Z(n15655)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i11996_2_lut_3_lut_4_lut.init = 16'hfff1;
    LUT4 i1850_1_lut_rep_422_2_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .Z(lastAddress_31__N_1310)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i1850_1_lut_rep_422_2_lut.init = 16'h1111;
    LUT4 lastAddress_i1_i22_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(lastAddress[21]), .D(SRAM_WE_N_1254), .Z(n43)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i22_3_lut_3_lut_4_lut.init = 16'hf011;
    CCU2D sub_991_add_2_11 (.A0(currPWMCount[9]), .B0(currPWMCountMax[9]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[10]), .B1(currPWMCountMax[10]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14078), .COUT(n14079));
    defparam sub_991_add_2_11.INIT0 = 16'h5999;
    defparam sub_991_add_2_11.INIT1 = 16'h5999;
    defparam sub_991_add_2_11.INJECT1_0 = "NO";
    defparam sub_991_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_991_add_2_9 (.A0(currPWMCount[7]), .B0(currPWMCountMax[7]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[8]), .B1(currPWMCountMax[8]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14077), .COUT(n14078));
    defparam sub_991_add_2_9.INIT0 = 16'h5999;
    defparam sub_991_add_2_9.INIT1 = 16'h5999;
    defparam sub_991_add_2_9.INJECT1_0 = "NO";
    defparam sub_991_add_2_9.INJECT1_1 = "NO";
    LUT4 lastAddress_i1_i32_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(lastAddress[31]), .D(SRAM_WE_N_1254), .Z(n33)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i32_3_lut_3_lut_4_lut.init = 16'hf011;
    CCU2D sub_991_add_2_7 (.A0(currPWMCount[5]), .B0(currPWMCountMax[5]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[6]), .B1(currPWMCountMax[6]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14076), .COUT(n14077));
    defparam sub_991_add_2_7.INIT0 = 16'h5999;
    defparam sub_991_add_2_7.INIT1 = 16'h5999;
    defparam sub_991_add_2_7.INJECT1_0 = "NO";
    defparam sub_991_add_2_7.INJECT1_1 = "NO";
    LUT4 lastAddress_i1_i24_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(lastAddress[23]), .D(SRAM_WE_N_1254), .Z(n41)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i24_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 lastAddress_i1_i23_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(lastAddress[22]), .D(SRAM_WE_N_1254), .Z(n42)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i23_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 lastAddress_i1_i30_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(lastAddress[29]), .D(SRAM_WE_N_1254), .Z(n35)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i30_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 lastAddress_i1_i29_3_lut_3_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(lastAddress[28]), .D(SRAM_WE_N_1254), .Z(n36)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam lastAddress_i1_i29_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i3346_2_lut_rep_364_3_lut_4_lut_3_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL_adj_2610[18]), .Z(BUS_ADDR_INTERNAL_18_derived_1)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[2] 137[9])
    defparam i3346_2_lut_rep_364_3_lut_4_lut_3_lut.init = 16'h5151;
    VLO i1 (.Z(GND_net));
    CCU2D sub_991_add_2_5 (.A0(currPWMCount[3]), .B0(currPWMCountMax[3]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[4]), .B1(currPWMCountMax[4]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14075), .COUT(n14076));
    defparam sub_991_add_2_5.INIT0 = 16'h5999;
    defparam sub_991_add_2_5.INIT1 = 16'h5999;
    defparam sub_991_add_2_5.INJECT1_0 = "NO";
    defparam sub_991_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(BUS_ADDR_INTERNAL_adj_2610[15]), .B(n18271), 
         .C(n17457), .D(BUS_addr[10]), .Z(n9)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i1_2_lut_4_lut.init = 16'hceff;
    LUT4 i10580_2_lut_4_lut (.A(BUS_ADDR_INTERNAL_adj_2610[15]), .B(n18271), 
         .C(n17457), .D(n17362), .Z(n13936)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i10580_2_lut_4_lut.init = 16'hce00;
    CCU2D sub_991_add_2_3 (.A0(currPWMCount[1]), .B0(currPWMCountMax[1]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[2]), .B1(currPWMCountMax[2]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14074), .COUT(n14075));
    defparam sub_991_add_2_3.INIT0 = 16'h5999;
    defparam sub_991_add_2_3.INIT1 = 16'h5999;
    defparam sub_991_add_2_3.INJECT1_0 = "NO";
    defparam sub_991_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_991_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(currPWMCount[0]), .B1(currPWMCountMax[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n14074));
    defparam sub_991_add_2_1.INIT0 = 16'h0000;
    defparam sub_991_add_2_1.INIT1 = 16'h5999;
    defparam sub_991_add_2_1.INJECT1_0 = "NO";
    defparam sub_991_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_675 (.A(BUS_DATA_INTERNAL_adj_2601[8]), .B(MDM_data[8]), 
         .C(n17330), .D(PIC_data[8]), .Z(BUS_data[8])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i2_4_lut_adj_675.init = 16'hffec;
    LUT4 i1_4_lut (.A(otherData[9]), .B(writeData[9]), .C(n17272), .D(n18278), 
         .Z(n4_adj_2532)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut.init = 16'hce0a;
    LUT4 i12105_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4265), .D(n4249), 
         .Z(n15767)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12105_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12601_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4616), .D(n4600), 
         .Z(n16263)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12601_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6863_2_lut (.A(BUS_req[2]), .B(BUS_currGrantID_3__N_74[0]), .Z(BUS_currGrantID_3__N_74[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(125[4] 131[11])
    defparam i6863_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_676 (.A(Sprite_readData2[10]), .B(writeData[10]), 
         .C(n14584), .D(n18278), .Z(n4_adj_2523)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_676.init = 16'hce0a;
    LUT4 i1_4_lut_adj_677 (.A(Sprite_readData2[11]), .B(writeData[11]), 
         .C(n14584), .D(n18278), .Z(n4)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_677.init = 16'hce0a;
    LUT4 i12600_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4581), .D(n4565), 
         .Z(n16262)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12600_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12598_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4615), .D(n4599), 
         .Z(n16260)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12598_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_336_4_lut (.A(BUS_ADDR_INTERNAL_adj_2610[16]), .B(n18277), 
         .C(n17457), .D(n17381), .Z(n17344)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i1_2_lut_rep_336_4_lut.init = 16'hffce;
    LUT4 i1_2_lut_rep_290_4_lut (.A(n15539), .B(n17458), .C(n17311), .D(n17373), 
         .Z(n17298)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i1_2_lut_rep_290_4_lut.init = 16'hfffb;
    LUT4 i2_3_lut_rep_297 (.A(n15534), .B(n17378), .C(n17376), .Z(n17305)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i2_3_lut_rep_297.init = 16'hfefe;
    LUT4 i13114_2_lut_4_lut (.A(n15534), .B(n17378), .C(n17376), .D(n18260), 
         .Z(n16497)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i13114_2_lut_4_lut.init = 16'h0001;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i7_4_lut (.A(n9), .B(n14_adj_2564), .C(n17411), .D(n17344), 
         .Z(n15534)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i7_4_lut.init = 16'hffef;
    LUT4 i6_4_lut (.A(n17377), .B(n17383), .C(n17379), .D(BUS_addr[11]), 
         .Z(n14_adj_2564)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_678 (.A(Sprite_readData2[12]), .B(writeData[12]), 
         .C(n14584), .D(n18278), .Z(n4_adj_2560)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_678.init = 16'hce0a;
    LUT4 i1_4_lut_adj_679 (.A(Sprite_readData2[13]), .B(writeData[13]), 
         .C(n14584), .D(n18278), .Z(n4_adj_2559)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_679.init = 16'hce0a;
    LUT4 i1_4_lut_adj_680 (.A(Sprite_readData2[14]), .B(writeData[14]), 
         .C(n14584), .D(n18278), .Z(n4_adj_2558)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_680.init = 16'hce0a;
    LUT4 i1_4_lut_adj_681 (.A(Sprite_readData2[15]), .B(writeData[15]), 
         .C(n14584), .D(n18278), .Z(n4_adj_2527)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_681.init = 16'hce0a;
    LUT4 i12597_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4580), .D(n4564), 
         .Z(n16259)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12597_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_4_lut_adj_682 (.A(BUS_DATA_INTERNAL_adj_2580[4]), .B(writeData[4]), 
         .C(n17274), .D(n18278), .Z(n4_adj_2568)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_682.init = 16'heca0;
    LUT4 i12595_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4614), .D(n4598), 
         .Z(n16257)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12595_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12573_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4609), .D(n4593), 
         .Z(n16235)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12573_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6894_2_lut_rep_317_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[9]), .D(BUS_ADDR_INTERNAL_adj_2610[9]), .Z(n17325)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6894_2_lut_rep_317_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i12106_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4300), .D(n4284), 
         .Z(n15768)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12106_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_302_3_lut_4_lut (.A(n18259), .B(n17423), .C(n17458), 
         .D(n17385), .Z(n17310)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i1_2_lut_rep_302_3_lut_4_lut.init = 16'hffef;
    LUT4 i7007_2_lut_3_lut_4_lut (.A(n18259), .B(n17423), .C(n17458), 
         .D(n17385), .Z(Sprite_pointers_N_1136)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i7007_2_lut_3_lut_4_lut.init = 16'hef0f;
    LUT4 i3_4_lut_adj_683 (.A(n5_adj_2567), .B(BUS_DATA_INTERNAL_adj_2601[1]), 
         .C(n161), .D(n17330), .Z(BUS_data[1])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i3_4_lut_adj_683.init = 16'hfefa;
    LUT4 i1_4_lut_adj_684 (.A(BUS_DATA_INTERNAL_adj_2609[1]), .B(n17274), 
         .C(OUT_ENABLE), .D(BUS_DATA_INTERNAL_adj_2580[1]), .Z(n5_adj_2567)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_684.init = 16'heca0;
    LUT4 i3_4_lut_adj_685 (.A(n5), .B(BUS_DATA_INTERNAL_adj_2601[2]), .C(n160), 
         .D(n17330), .Z(BUS_data[2])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i3_4_lut_adj_685.init = 16'hfefa;
    LUT4 i1_4_lut_adj_686 (.A(BUS_DATA_INTERNAL_adj_2609[2]), .B(n17274), 
         .C(OUT_ENABLE), .D(BUS_DATA_INTERNAL_adj_2580[2]), .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_686.init = 16'heca0;
    LUT4 BUS_ADDR_IN_1__I_0_805_i3_2_lut_rep_304_3_lut_3_lut_4_lut (.A(n18259), 
         .B(n17423), .C(n17458), .D(n17385), .Z(n17312)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam BUS_ADDR_IN_1__I_0_805_i3_2_lut_rep_304_3_lut_3_lut_4_lut.init = 16'hefff;
    LUT4 i3_4_lut_adj_687 (.A(n5_adj_2563), .B(BUS_DATA_INTERNAL_adj_2601[3]), 
         .C(n159), .D(n17330), .Z(BUS_data[3])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i3_4_lut_adj_687.init = 16'hfefa;
    LUT4 i1_4_lut_adj_688 (.A(BUS_DATA_INTERNAL_adj_2609[3]), .B(n17274), 
         .C(OUT_ENABLE), .D(BUS_DATA_INTERNAL_adj_2580[3]), .Z(n5_adj_2563)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_688.init = 16'heca0;
    LUT4 i1_4_lut_adj_689 (.A(BUS_DATA_INTERNAL_adj_2580[5]), .B(writeData[5]), 
         .C(n17274), .D(n18278), .Z(n4_adj_2524)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_689.init = 16'heca0;
    LUT4 i1_4_lut_adj_690 (.A(BUS_DATA_INTERNAL_adj_2580[6]), .B(writeData[6]), 
         .C(n17274), .D(n18278), .Z(n4_adj_2565)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_690.init = 16'heca0;
    LUT4 i1_4_lut_adj_691 (.A(BUS_DATA_INTERNAL_adj_2580[7]), .B(writeData[7]), 
         .C(n17274), .D(n18278), .Z(n4_adj_2562)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(104[14:49])
    defparam i1_4_lut_adj_691.init = 16'heca0;
    LUT4 BUS_ADDR_IN_1__I_0_807_i3_2_lut_rep_294_2_lut_3_lut_3_lut_4_lut (.A(n18259), 
         .B(n17423), .C(n17458), .D(n17385), .Z(n17302)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam BUS_ADDR_IN_1__I_0_807_i3_2_lut_rep_294_2_lut_3_lut_3_lut_4_lut.init = 16'hff1f;
    LUT4 i2_2_lut_3_lut_3_lut_2_lut_3_lut_3_lut_4_lut (.A(n18259), .B(n17423), 
         .C(n17458), .D(n17385), .Z(n10346)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[15:23])
    defparam i2_2_lut_3_lut_3_lut_2_lut_3_lut_3_lut_4_lut.init = 16'hef1f;
    LUT4 lastAddress_i1_i16_3_lut_4_lut (.A(n17355), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[15]), .Z(n49)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i16_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i12675_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4371), .D(n4355), 
         .Z(n16337)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12675_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12641_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4476), .D(n4460), 
         .Z(n16303)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12641_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12642_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4511), .D(n4495), 
         .Z(n16304)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12642_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12604_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4503), .D(n4487), 
         .Z(n16266)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12604_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12603_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4468), .D(n4452), 
         .Z(n16265)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12603_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12676_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4406), .D(n4390), 
         .Z(n16338)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12676_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12679_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4293), .D(n4277), 
         .Z(n16341)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12679_3_lut_4_lut.init = 16'hf4b0;
    LUT4 lastAddress_i1_i7_3_lut_4_lut (.A(n17374), .B(n17458), .C(SRAM_WE_N_1254), 
         .D(lastAddress[6]), .Z(n58)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam lastAddress_i1_i7_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i12678_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4258), .D(n4242), 
         .Z(n16340)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12678_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12673_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4405), .D(n4389), 
         .Z(n16335)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12673_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12672_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4370), .D(n4354), 
         .Z(n16334)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12672_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12670_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4404), .D(n4388), 
         .Z(n16332)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12670_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12669_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4369), .D(n4353), 
         .Z(n16331)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12669_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i2_4_lut_4_lut_4_lut_adj_692 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[10]), .D(BUS_ADDR_INTERNAL_adj_2610[10]), 
         .Z(BUS_addr[10])) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i2_4_lut_4_lut_4_lut_adj_692.init = 16'h7531;
    LUT4 i12667_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4403), .D(n4387), 
         .Z(n16329)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12667_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12666_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4368), .D(n4352), 
         .Z(n16328)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12666_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12664_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4402), .D(n4386), 
         .Z(n16326)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12664_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_currGrantID_1__I_0_i3_4_lut (.A(BUS_currGrantID_3__N_74[0]), 
         .B(BUS_req[2]), .C(BUS_currGrantID[1]), .D(BUS_currGrantID[0]), 
         .Z(BUS_currGrantID_3__N_55)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (B (D)+!B (C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(119[13:50])
    defparam BUS_currGrantID_1__I_0_i3_4_lut.init = 16'hf530;
    LUT4 i12663_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4367), .D(n4351), 
         .Z(n16325)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12663_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12654_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4401), .D(n4385), 
         .Z(n16316)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12654_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12653_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4366), .D(n4350), 
         .Z(n16315)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12653_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12651_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4400), .D(n4384), 
         .Z(n16313)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12651_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12650_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4365), .D(n4349), 
         .Z(n16312)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12650_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12648_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4399), .D(n4383), 
         .Z(n16310)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12648_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12647_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4364), .D(n4348), 
         .Z(n16309)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12647_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12645_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4398), .D(n4382), 
         .Z(n16307)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12645_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12644_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4363), .D(n4347), 
         .Z(n16306)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12644_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12632_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4510), .D(n4494), 
         .Z(n16294)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12632_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12631_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4475), .D(n4459), 
         .Z(n16293)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12631_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12629_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4509), .D(n4493), 
         .Z(n16291)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12629_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12628_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4474), .D(n4458), 
         .Z(n16290)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12628_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12626_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4508), .D(n4492), 
         .Z(n16288)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12626_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12625_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4473), .D(n4457), 
         .Z(n16287)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12625_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12623_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4507), .D(n4491), 
         .Z(n16285)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12623_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12622_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4472), .D(n4456), 
         .Z(n16284)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12622_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12620_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4506), .D(n4490), 
         .Z(n16282)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12620_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12619_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4471), .D(n4455), 
         .Z(n16281)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12619_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12617_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4505), .D(n4489), 
         .Z(n16279)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12617_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12616_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4470), .D(n4454), 
         .Z(n16278)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12616_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12614_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4504), .D(n4488), 
         .Z(n16276)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12614_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i11976_2_lut (.A(currPixel[2]), .B(currPixel[4]), .Z(n15633)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11976_2_lut.init = 16'heeee;
    PLL PLL_Ent (.LOGIC_CLOCK_N_57(LOGIC_CLOCK_N_57), .LOGIC_CLOCK(LOGIC_CLOCK), 
        .CLK_c(CLK_c), .PIXEL_CLOCK(PIXEL_CLOCK), .GND_net(GND_net), .PIXEL_CLOCK_N_293(PIXEL_CLOCK_N_293)) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(244[10:13])
    LUT4 i12613_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4469), .D(n4453), 
         .Z(n16275)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12613_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12594_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4579), .D(n4563), 
         .Z(n16256)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12594_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12585_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4613), .D(n4597), 
         .Z(n16247)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12585_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12584_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4578), .D(n4562), 
         .Z(n16246)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12584_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12582_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4612), .D(n4596), 
         .Z(n16244)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12582_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12581_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4577), .D(n4561), 
         .Z(n16243)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12581_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12579_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4611), .D(n4595), 
         .Z(n16241)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12579_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12578_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4576), .D(n4560), 
         .Z(n16240)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12578_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12576_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4610), .D(n4594), 
         .Z(n16238)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12576_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i6795_2_lut_3_lut_rep_473 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[10]), .Z(n18269)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(99[26:48])
    defparam i6795_2_lut_3_lut_rep_473.init = 16'h2020;
    LUT4 i12575_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4575), .D(n4559), 
         .Z(n16237)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12575_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12109_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4301), .D(n4285), 
         .Z(n15771)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12109_3_lut_4_lut.init = 16'hf4b0;
    MatrixBusHandler MDM (.VRAM_DATA_OUT({VRAM_DATA_OUT}), .GND_net(GND_net), 
            .LOGIC_CLOCK(LOGIC_CLOCK), .n17458(n17458), .n17411(n17411), 
            .n18270(n18270), .n17382(n17382), .lastAddress_31__N_1338(lastAddress_31__N_1338), 
            .\BUS_DATA_INTERNAL[7] (BUS_DATA_INTERNAL_adj_2580[7]), .yOffset({Open_75, 
            Open_76, Open_77, Open_78, Open_79, Open_80, Open_81, 
            yOffset[0]}), .n17339(n17339), .n17333(n17333), .n17332(n17332), 
            .n17331(n17331), .BUS_data({BUS_data}), .n4305(n4305), .n4306(n4306), 
            .n4307(n4307), .n4308(n4308), .\state[0] (state[0]), .\BUS_DATA_INTERNAL[6] (BUS_DATA_INTERNAL_adj_2580[6]), 
            .n17276(n17276), .n17314(n17314), .n17334(n17334), .n17321(n17321), 
            .n17312(n17312), .\BUS_DATA_INTERNAL[5] (BUS_DATA_INTERNAL_adj_2580[5]), 
            .\SpriteRead_yInSprite_7__N_597[0] (SpriteRead_yInSprite_7__N_597[0]), 
            .\VRAM_ADDR[0] (VRAM_ADDR[0]), .\BUS_DATA_INTERNAL[4] (BUS_DATA_INTERNAL_adj_2580[4]), 
            .n4608(n4608), .n4609(n4609), .n4610(n4610), .n4611(n4611), 
            .n4612(n4612), .n4613(n4613), .n4614(n4614), .n4615(n4615), 
            .n4616(n4616), .n4617(n4617), .n4618(n4618), .n4619(n4619), 
            .n4573(n4573), .n4574(n4574), .n4575(n4575), .n4576(n4576), 
            .n4591(n4591), .n17381(n17381), .lastAddress_31__N_1323(lastAddress_31__N_1323), 
            .n4577(n4577), .n4578(n4578), .n4579(n4579), .n4580(n4580), 
            .n4581(n4581), .n4582(n4582), .n4583(n4583), .n4584(n4584), 
            .n4592(n4592), .n4593(n4593), .n4594(n4594), .n4595(n4595), 
            .n4625(n4625), .n4596(n4596), .n4597(n4597), .n4598(n4598), 
            .n4599(n4599), .n4600(n4600), .n4601(n4601), .n4602(n4602), 
            .n4603(n4603), .n2877(n2877), .\BUS_DATA_INTERNAL[3] (BUS_DATA_INTERNAL_adj_2580[3]), 
            .n4557(n4557), .n4558(n4558), .n4559(n4559), .n4560(n4560), 
            .n4590(n4590), .n4561(n4561), .n4562(n4562), .n4563(n4563), 
            .n4564(n4564), .n17373(n17373), .lastAddress_31__N_1413(lastAddress_31__N_1413), 
            .n2878(n2878), .\BUS_DATA_INTERNAL[2] (BUS_DATA_INTERNAL_adj_2580[2]), 
            .n2879(n2879), .\BUS_DATA_INTERNAL[1] (BUS_DATA_INTERNAL_adj_2580[1]), 
            .SpriteRead_yValid_N_1158({Open_82, Open_83, Open_84, Open_85, 
            SpriteRead_yValid_N_1158[3:2], Open_86, Open_87}), .n2880(n2880), 
            .\BUS_DATA_INTERNAL[0] (BUS_DATA_INTERNAL_adj_2580[0]), .n4604(n4604), 
            .n4605(n4605), .n4606(n4606), .n4607(n4607), .VRAM_WC(VRAM_WC), 
            .n8(n8), .VRAM_DATA({VRAM_DATA}), .\BUS_ADDR_INTERNAL[0] (BUS_ADDR_INTERNAL[0]), 
            .n4355(n4355), .n4356(n4356), .n4357(n4357), .n4358(n4358), 
            .n4460(n4460), .n4461(n4461), .n4462(n4462), .n4463(n4463), 
            .n4565(n4565), .n4566(n4566), .n4567(n4567), .n4568(n4568), 
            .Sprite_pointers_N_1123(Sprite_pointers_N_1123), .VCC_net(VCC_net), 
            .n4250(n4250), .n4251(n4251), .n4252(n4252), .n4253(n4253), 
            .n17342(n17342), .n17310(n17310), .n4569(n4569), .n4570(n4570), 
            .n4571(n4571), .n4572(n4572), .n4585(n4585), .n4586(n4586), 
            .n4587(n4587), .n4588(n4588), .n4620(n4620), .n4621(n4621), 
            .n4622(n4622), .n4623(n4623), .n4503(n4503), .n4504(n4504), 
            .n4505(n4505), .n4506(n4506), .\Sprite_readData2[10] (Sprite_readData2[10]), 
            .n4507(n4507), .n4508(n4508), .n4509(n4509), .n4510(n4510), 
            .n17371(n17371), .lastAddress_31__N_1337(lastAddress_31__N_1337), 
            .\Sprite_readData2[11] (Sprite_readData2[11]), .\Sprite_readData2[12] (Sprite_readData2[12]), 
            .\Sprite_readData2[13] (Sprite_readData2[13]), .n4511(n4511), 
            .n4512(n4512), .n4513(n4513), .n4514(n4514), .n4468(n4468), 
            .n4469(n4469), .n4470(n4470), .n4471(n4471), .n4472(n4472), 
            .n4473(n4473), .n4474(n4474), .n4475(n4475), .n4476(n4476), 
            .n4477(n4477), .n4478(n4478), .n4479(n4479), .n18280(n18280), 
            .\Sprite_readData2[14] (Sprite_readData2[14]), .\Sprite_readData2[15] (Sprite_readData2[15]), 
            .latchMode({latchMode}), .n17343(n17343), .n4487(n4487), .n4488(n4488), 
            .n4489(n4489), .n4490(n4490), .xOffset({Open_88, Open_89, 
            Open_90, Open_91, Open_92, Open_93, xOffset[1:0]}), .VRAM_WE(VRAM_WE), 
            .\state[1] (state[1]), .n4491(n4491), .n4492(n4492), .n4493(n4493), 
            .n4494(n4494), .n4495(n4495), .n4496(n4496), .n4497(n4497), 
            .n4498(n4498), .n4452(n4452), .n4453(n4453), .n4454(n4454), 
            .n4455(n4455), .n17366(n17366), .MATRIX_CURRROW({MATRIX_CURRROW}), 
            .\BUS_ADDR_INTERNAL[3] (BUS_ADDR_INTERNAL_adj_2610[3]), .\BUS_currGrantID[0] (BUS_currGrantID[0]), 
            .\BUS_currGrantID[1] (BUS_currGrantID[1]), .\BUS_ADDR_INTERNAL[3]_adj_2 (BUS_ADDR_INTERNAL[3]), 
            .n17453(n17453), .n17326(n17326), .\BUS_ADDR_INTERNAL[14] (BUS_ADDR_INTERNAL[14]), 
            .\BUS_ADDR_INTERNAL[14]_adj_3 (BUS_ADDR_INTERNAL_adj_2610[14]), 
            .n17383(n17383), .\BUS_ADDR_INTERNAL[2] (BUS_ADDR_INTERNAL[2]), 
            .\BUS_ADDR_INTERNAL[2]_adj_4 (BUS_ADDR_INTERNAL_adj_2610[2]), 
            .\BUS_ADDR_INTERNAL[17] (BUS_ADDR_INTERNAL[17]), .\BUS_ADDR_INTERNAL[17]_adj_5 (BUS_ADDR_INTERNAL_adj_2610[17]), 
            .n18260(n18260), .n17272(n17272), .\BUS_ADDR_INTERNAL[5] (BUS_ADDR_INTERNAL[5]), 
            .\BUS_ADDR_INTERNAL[5]_adj_6 (BUS_ADDR_INTERNAL_adj_2610[5]), 
            .n17380(n17380), .n4456(n4456), .n4457(n4457), .n4458(n4458), 
            .n4459(n4459), .\BUS_ADDR_INTERNAL[13] (BUS_ADDR_INTERNAL[13]), 
            .\BUS_ADDR_INTERNAL[13]_adj_7 (BUS_ADDR_INTERNAL_adj_2610[13]), 
            .n17379(n17379), .\BUS_ADDR_INTERNAL[8] (BUS_ADDR_INTERNAL[8]), 
            .\BUS_ADDR_INTERNAL[8]_adj_8 (BUS_ADDR_INTERNAL_adj_2610[8]), 
            .n17378(n17378), .\BUS_ADDR_INTERNAL[9] (BUS_ADDR_INTERNAL[9]), 
            .\BUS_ADDR_INTERNAL[9]_adj_9 (BUS_ADDR_INTERNAL_adj_2610[9]), 
            .n17376(n17376), .\BUS_ADDR_INTERNAL[4] (BUS_ADDR_INTERNAL[4]), 
            .\BUS_ADDR_INTERNAL[4]_adj_10 (BUS_ADDR_INTERNAL_adj_2610[4]), 
            .n17375(n17375), .n17275(n17275), .\state[1]_adj_11 (state_adj_2613[1]), 
            .n17434(n17434), .n17457(n17457), .n15469(n15469), .\BUS_ADDR_INTERNAL[6] (BUS_ADDR_INTERNAL[6]), 
            .\BUS_ADDR_INTERNAL[6]_adj_12 (BUS_ADDR_INTERNAL_adj_2610[6]), 
            .n17374(n17374), .\BUS_ADDR_INTERNAL[7] (BUS_ADDR_INTERNAL[7]), 
            .\BUS_ADDR_INTERNAL[7]_adj_13 (BUS_ADDR_INTERNAL_adj_2610[7]), 
            .\BUS_ADDR_INTERNAL[12] (BUS_ADDR_INTERNAL[12]), .\BUS_ADDR_INTERNAL[12]_adj_14 (BUS_ADDR_INTERNAL_adj_2610[12]), 
            .n17377(n17377), .n17407(n17407), .\BUS_ADDR_INTERNAL[16] (BUS_ADDR_INTERNAL[16]), 
            .\BUS_ADDR_INTERNAL[16]_adj_15 (BUS_ADDR_INTERNAL_adj_2610[16]), 
            .n17362(n17362), .\BUS_ADDR_INTERNAL[15] (BUS_ADDR_INTERNAL[15]), 
            .\BUS_ADDR_INTERNAL[15]_adj_16 (BUS_ADDR_INTERNAL_adj_2610[15]), 
            .n17355(n17355), .\state[3] (state[3]), .\yOffset[3] (yOffset[3]), 
            .\yOffset[2] (yOffset[2]), .\yOffset[1] (yOffset[1]), .n16084(n16084), 
            .n16085(n16085), .n4499(n4499), .n4500(n4500), .n4501(n4501), 
            .n4502(n4502), .n16097(n16097), .n16098(n16098), .n16107(n16107), 
            .n16108(n16108), .n33(n33_adj_2561), .\BUS_ADDR_INTERNAL[0]_adj_17 (BUS_ADDR_INTERNAL_adj_2610[0]), 
            .n17385(n17385), .n16114(n16114), .n16115(n16115), .n4464(n4464), 
            .n4465(n4465), .n4466(n4466), .n4467(n4467), .n4480(n4480), 
            .n4481(n4481), .n4482(n4482), .n4483(n4483), .n4515(n4515), 
            .n4516(n4516), .n4517(n4517), .n4518(n4518), .n9891(n9891), 
            .n4398(n4398), .n4399(n4399), .n4400(n4400), .n4401(n4401), 
            .BUS_DONE_OUT_N_1051(BUS_DONE_OUT_N_1051), .n4402(n4402), .n4403(n4403), 
            .n4404(n4404), .n4405(n4405), .n4406(n4406), .n4407(n4407), 
            .n4408(n4408), .n4409(n4409), .n4363(n4363), .n4364(n4364), 
            .n4365(n4365), .n4366(n4366), .n4367(n4367), .n4368(n4368), 
            .n4369(n4369), .n4370(n4370), .n4371(n4371), .n4372(n4372), 
            .n4373(n4373), .n4374(n4374), .n4382(n4382), .n4383(n4383), 
            .n4384(n4384), .n4385(n4385), .n4386(n4386), .n4387(n4387), 
            .n4388(n4388), .n4389(n4389), .n16121(n16121), .n16122(n16122), 
            .n4390(n4390), .n4391(n4391), .n4392(n4392), .n4393(n4393), 
            .n4347(n4347), .n4348(n4348), .n4349(n4349), .n4350(n4350), 
            .n4351(n4351), .n4352(n4352), .n4353(n4353), .n4354(n4354), 
            .n16126(n16126), .n16127(n16127), .n16128(n16128), .n16129(n16129), 
            .n16130(n16130), .n16131(n16131), .n4394(n4394), .n4395(n4395), 
            .n4396(n4396), .n4397(n4397), .n16132(n16132), .n16133(n16133), 
            .n4359(n4359), .n4360(n4360), .n4361(n4361), .n4362(n4362), 
            .n4375(n4375), .n4376(n4376), .n4377(n4377), .n4378(n4378), 
            .n17329(n17329), .n17327(n17327), .n16141(n16141), .n16142(n16142), 
            .n4410(n4410), .n4411(n4411), .n4412(n4412), .n4413(n4413), 
            .n4293(n4293), .n4294(n4294), .n4295(n4295), .n4296(n4296), 
            .n4297(n4297), .n4298(n4298), .n4299(n4299), .n4300(n4300), 
            .n4301(n4301), .n4302(n4302), .n4303(n4303), .n4304(n4304), 
            .n4258(n4258), .n4259(n4259), .n4260(n4260), .n4261(n4261), 
            .n4262(n4262), .n4263(n4263), .n4264(n4264), .n4265(n4265), 
            .n4266(n4266), .n4267(n4267), .n4268(n4268), .n4269(n4269), 
            .n4277(n4277), .n4278(n4278), .n4279(n4279), .n4280(n4280), 
            .n4281(n4281), .n4282(n4282), .n4283(n4283), .n4284(n4284), 
            .n4285(n4285), .n4286(n4286), .n4287(n4287), .n4288(n4288), 
            .n4242(n4242), .n4243(n4243), .n4244(n4244), .n4245(n4245), 
            .n4246(n4246), .n4247(n4247), .n4248(n4248), .n4249(n4249), 
            .n17279(n17279), .n17274(n17274), .n16143(n16143), .n16144(n16144), 
            .n4289(n4289), .n4290(n4290), .n4291(n4291), .n4292(n4292), 
            .n16145(n16145), .n16146(n16146), .n4254(n4254), .n4255(n4255), 
            .n4256(n4256), .n4257(n4257), .n4270(n4270), .n4271(n4271), 
            .n4272(n4272), .n4273(n4273), .n16147(n16147), .n16148(n16148), 
            .n16156(n16156), .n16157(n16157), .Sprite_pointers_N_1136(Sprite_pointers_N_1136), 
            .n17287(n17287), .n16158(n16158), .n16159(n16159), .SpriteRead_yInSprite({SpriteRead_yInSprite}), 
            .LOGIC_CLOCK_enable_52(LOGIC_CLOCK_enable_52), .\SpriteRead_yValid_N_1158[1] (SpriteRead_yValid_N_1158[1]), 
            .n16160(n16160), .n16161(n16161), .n16162(n16162), .n16163(n16163), 
            .n16171(n16171), .n16172(n16172), .n18264(n18264), .\BUS_ADDR_INTERNAL[18] (BUS_ADDR_INTERNAL_adj_2610[18]), 
            .lastAddress_31__N_1310(lastAddress_31__N_1310), .n18271(n18271), 
            .n18277(n18277), .n18266(n18266), .n18262(n18262), .n16173(n16173), 
            .n16174(n16174), .n16175(n16175), .n16176(n16176), .\BUS_ADDR_INTERNAL[11] (BUS_ADDR_INTERNAL_adj_2610[11]), 
            .n18273(n18273), .n18272(n18272), .n16177(n16177), .n16178(n16178), 
            .n18268(n18268), .\BUS_ADDR_INTERNAL[10] (BUS_ADDR_INTERNAL_adj_2610[10]), 
            .n18269(n18269), .n18267(n18267), .n15749(n15749), .n15750(n15750), 
            .n16186(n16186), .n16187(n16187), .n16188(n16188), .n16189(n16189), 
            .n16190(n16190), .n16191(n16191), .\BUS_currGrantID_3__N_74[0] (BUS_currGrantID_3__N_74[0]), 
            .n17408(n17408), .n17368(n17368), .n16192(n16192), .n16193(n16193), 
            .n17452(n17452), .n16201(n16201), .n16202(n16202), .n16203(n16203), 
            .n16204(n16204), .n16205(n16205), .n16206(n16206), .n16207(n16207), 
            .n16208(n16208), .\BUS_ADDR_INTERNAL[18]_derived_1 (BUS_ADDR_INTERNAL_18_derived_1), 
            .n2504(n2504), .n15752(n15752), .n15753(n15753), .lastAddress_31__N_1425(lastAddress_31__N_1425), 
            .n17384(n17384), .n6250(n6250), .n17311(n17311), .n15755(n15755), 
            .n15756(n15756), .n15758(n15758), .n15759(n15759), .n15761(n15761), 
            .n15762(n15762), .n16216(n16216), .n16217(n16217), .n16218(n16218), 
            .n16219(n16219), .n16220(n16220), .n16221(n16221), .n16222(n16222), 
            .n16223(n16223), .reset(reset), .state_7__N_345(state_7__N_345), 
            .\Sprite_readAddr_13__N_752[13] (Sprite_readAddr_13__N_752[13]), 
            .n17313(n17313), .\Sprite_readAddr_13__N_752[11] (Sprite_readAddr_13__N_752[11]), 
            .\Sprite_readAddr_13__N_752[12] (Sprite_readAddr_13__N_752[12]), 
            .\Sprite_readAddr_13__N_752[9] (Sprite_readAddr_13__N_752[9]), 
            .\Sprite_readAddr_13__N_752[10] (Sprite_readAddr_13__N_752[10]), 
            .n15764(n15764), .n15765(n15765), .n16231(n16231), .n16232(n16232), 
            .n16234(n16234), .n16235(n16235), .\Sprite_readAddr_13__N_752[7] (Sprite_readAddr_13__N_752[7]), 
            .\Sprite_readAddr_13__N_752[8] (Sprite_readAddr_13__N_752[8]), 
            .\Sprite_readAddr_13__N_752[5] (Sprite_readAddr_13__N_752[5]), 
            .\Sprite_readAddr_13__N_752[6] (Sprite_readAddr_13__N_752[6]), 
            .\Sprite_readAddr_13__N_752[3] (Sprite_readAddr_13__N_752[3]), 
            .\Sprite_readAddr_13__N_752[4] (Sprite_readAddr_13__N_752[4]), 
            .\Sprite_readAddr_13__N_752[1] (Sprite_readAddr_13__N_752[1]), 
            .\Sprite_readAddr_13__N_752[2] (Sprite_readAddr_13__N_752[2]), 
            .n16237(n16237), .n16238(n16238), .\Sprite_readAddr_13__N_752[0] (Sprite_readAddr_13__N_752[0]), 
            .n17256(n17256), .n16240(n16240), .n16241(n16241), .n16243(n16243), 
            .n16244(n16244), .n16246(n16246), .n16247(n16247), .n16251(n16251), 
            .n16252(n16252), .n16256(n16256), .n16257(n16257), .n16259(n16259), 
            .n16260(n16260), .n16262(n16262), .n16263(n16263), .n15767(n15767), 
            .n15768(n15768), .n16265(n16265), .n16266(n16266), .n15770(n15770), 
            .n15771(n15771), .n16270(n16270), .n16271(n16271), .n16275(n16275), 
            .n16276(n16276), .n16278(n16278), .n16279(n16279), .n16281(n16281), 
            .n16282(n16282), .\VRAM_ADDR[1] (VRAM_ADDR[1]), .\VRAM_ADDR[2] (VRAM_ADDR[2]), 
            .\VRAM_ADDR[3] (VRAM_ADDR[3]), .\VRAM_ADDR[4] (VRAM_ADDR[4]), 
            .\VRAM_ADDR[5] (VRAM_ADDR[5]), .\VRAM_ADDR[6] (VRAM_ADDR[6]), 
            .\VRAM_ADDR[7] (VRAM_ADDR[7]), .\VRAM_ADDR[8] (VRAM_ADDR[8]), 
            .\BUS_ADDR_INTERNAL[1] (BUS_ADDR_INTERNAL[1]), .\BUS_ADDR_INTERNAL[10]_adj_18 (BUS_ADDR_INTERNAL[10]), 
            .\BUS_ADDR_INTERNAL[11]_adj_19 (BUS_ADDR_INTERNAL[11]), .n16284(n16284), 
            .n16285(n16285), .n16287(n16287), .n16288(n16288), .n17337(n17337), 
            .n17325(n17325), .\BUS_addr[10] (BUS_addr[10]), .\BUS_addr[11] (BUS_addr[11]), 
            .n17335(n17335), .n17338(n17338), .\xOffset[2] (xOffset[2]), 
            .\xOffset[3] (xOffset[3]), .n9(n9_adj_2566), .n16290(n16290), 
            .n16291(n16291), .n17340(n17340), .n15655(n15655), .n16293(n16293), 
            .n16294(n16294), .n15436(n15436), .n2642(n2642), .n16298(n16298), 
            .n16299(n16299), .n16303(n16303), .n16304(n16304), .n16306(n16306), 
            .n16307(n16307), .n16309(n16309), .n16310(n16310), .n16312(n16312), 
            .n16313(n16313), .n16315(n16315), .n16316(n16316), .n16320(n16320), 
            .n16321(n16321), .n4(n4_adj_2525), .n17305(n17305), .n17298(n17298), 
            .n63(n63_adj_2556), .n63_adj_20(n63_adj_2557), .n16325(n16325), 
            .n16326(n16326), .n16328(n16328), .n16329(n16329), .n16331(n16331), 
            .n16332(n16332), .n16334(n16334), .n16335(n16335), .n16337(n16337), 
            .n16338(n16338), .lastAddress_31__N_1434(lastAddress_31__N_1434), 
            .n17302(n17302), .n17309(n17309), .n17308(n17308), .n16340(n16340), 
            .n16341(n16341), .\currSprite_size[6] (currSprite_size[6]), 
            .\currSprite_size[7] (currSprite_size[7]), .lastAddress_31__N_1401(lastAddress_31__N_1401), 
            .\currSprite_size[4] (currSprite_size[4]), .\currSprite_size[5] (currSprite_size[5]), 
            .lastAddress_31__N_1336(lastAddress_31__N_1336), .n17304(n17304), 
            .n7(n7), .n18276(n18276), .n18274(n18274), .\currSprite_size[2] (currSprite_size[2]), 
            .\currSprite_size[3] (currSprite_size[3]), .n18275(n18275), 
            .n18265(n18265), .n18263(n18263), .n17409(n17409), .n17423(n17423), 
            .n18259(n18259), .n17394(n17394), .\currSprite_size[1] (currSprite_size[1]), 
            .lastAddress_31__N_1422(lastAddress_31__N_1422), .\MDM_data[8] (MDM_data[8]), 
            .\otherData[9] (otherData[9]), .n15539(n15539), .n17328(n17328), 
            .n6340(n6340), .SRAM_WE_N_1254(SRAM_WE_N_1254), .\lastAddress[18] (lastAddress[18]), 
            .n46(n46), .lastAddress_31__N_1431(lastAddress_31__N_1431), 
            .lastAddress_31__N_1383(lastAddress_31__N_1383), .lastAddress_31__N_1325(lastAddress_31__N_1325), 
            .lastAddress_31__N_1334(lastAddress_31__N_1334), .lastAddress_31__N_1326(lastAddress_31__N_1326), 
            .lastAddress_31__N_1404(lastAddress_31__N_1404), .lastAddress_31__N_1333(lastAddress_31__N_1333), 
            .lastAddress_31__N_1335(lastAddress_31__N_1335), .lastAddress_31__N_1330(lastAddress_31__N_1330), 
            .lastAddress_31__N_1419(lastAddress_31__N_1419), .lastAddress_31__N_1407(lastAddress_31__N_1407), 
            .lastAddress_31__N_1395(lastAddress_31__N_1395), .lastAddress_31__N_1386(lastAddress_31__N_1386), 
            .lastAddress_31__N_1331(lastAddress_31__N_1331), .lastAddress_31__N_1389(lastAddress_31__N_1389), 
            .lastAddress_31__N_1398(lastAddress_31__N_1398), .lastAddress_31__N_1328(lastAddress_31__N_1328), 
            .lastAddress_31__N_1392(lastAddress_31__N_1392), .lastAddress_31__N_1327(lastAddress_31__N_1327), 
            .lastAddress_31__N_1428(lastAddress_31__N_1428), .lastAddress_31__N_1339(lastAddress_31__N_1339), 
            .lastAddress_31__N_1332(lastAddress_31__N_1332), .lastAddress_31__N_1329(lastAddress_31__N_1329), 
            .lastAddress_31__N_1324(lastAddress_31__N_1324), .lastAddress_31__N_1340(lastAddress_31__N_1340), 
            .lastAddress_31__N_1416(lastAddress_31__N_1416), .lastAddress_31__N_1410(lastAddress_31__N_1410), 
            .n14584(n14584), .\SpriteRead_yValid_N_1158[4] (SpriteRead_yValid_N_1158[4]), 
            .n17299(n17299), .n17307(n17307), .n15549(n15549), .\SpriteRead_yValid_N_1158[0] (SpriteRead_yValid_N_1158[0]), 
            .n15571(n15571), .n8_adj_21(n8_adj_2526), .WRITE_DONE(WRITE_DONE_adj_2554), 
            .n10346(n10346), .n17456(n17456), .n17344(n17344), .RED_WRITE({RED_WRITE}), 
            .GREEN_WRITE({GREEN_WRITE}), .LOGIC_CLOCK_N_57(LOGIC_CLOCK_N_57), 
            .n17387(n17387), .BLUE_WRITE({BLUE_WRITE}), .ALPHA_WRITE({ALPHA_WRITE}));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(172[7:35])
    PIC PIC_BUS_INTERFACE (.PIC_DATA_IN_out_7(PIC_DATA_IN_out_7), .\BUS_currGrantID[1] (BUS_currGrantID[1]), 
        .\BUS_currGrantID[0] (BUS_currGrantID[0]), .\BUS_ADDR_INTERNAL[11] (BUS_ADDR_INTERNAL_adj_2610[11]), 
        .n18273(n18273), .\BUS_ADDR_INTERNAL[12] (BUS_ADDR_INTERNAL_adj_2610[12]), 
        .n18272(n18272), .GND_net(GND_net), .writeData({writeData[15:11], 
        Open_94, Open_95, Open_96, Open_97, Open_98, Open_99, Open_100, 
        Open_101, Open_102, Open_103, Open_104}), .LOGIC_CLOCK(LOGIC_CLOCK), 
        .PIC_DATA_IN_out_15(PIC_DATA_IN_out_15), .PIC_DATA_IN_out_14(PIC_DATA_IN_out_14), 
        .PIC_DATA_IN_out_13(PIC_DATA_IN_out_13), .PIC_DATA_IN_out_12(PIC_DATA_IN_out_12), 
        .PIC_DATA_IN_out_11(PIC_DATA_IN_out_11), .\BUS_ADDR_INTERNAL[9] (BUS_ADDR_INTERNAL_adj_2610[9]), 
        .n18268(n18268), .\BUS_ADDR_INTERNAL[10] (BUS_ADDR_INTERNAL_adj_2610[10]), 
        .n18269(n18269), .\BUS_ADDR_INTERNAL[8] (BUS_ADDR_INTERNAL_adj_2610[8]), 
        .n18267(n18267), .OUT_ENABLE(OUT_ENABLE), .n9950(n9950), .\PIC_data[0] (PIC_data[0]), 
        .\writeData[10] (writeData[10]), .PIC_DATA_IN_out_10(PIC_DATA_IN_out_10), 
        .\writeData[9] (writeData[9]), .PIC_DATA_IN_out_9(PIC_DATA_IN_out_9), 
        .\writeData[8] (writeData[8]), .PIC_DATA_IN_out_8(PIC_DATA_IN_out_8), 
        .n17298(n17298), .n17337(n17337), .n17325(n17325), .n15534(n15534), 
        .state({Open_105, Open_106, Open_107, state_adj_2613[4], Open_108, 
        Open_109, state_adj_2613[1], Open_110}), .n17270(n17270), .PIC_WE_IN_c(PIC_WE_IN_c), 
        .\BUS_data[0] (BUS_data[0]), .\BUS_ADDR_INTERNAL[0] (BUS_ADDR_INTERNAL_adj_2610[0]), 
        .PIC_ADDR_IN_c_0(PIC_ADDR_IN_c_0), .\BUS_ADDR_INTERNAL[1] (BUS_ADDR_INTERNAL_adj_2610[1]), 
        .\BUS_ADDR_INTERNAL[1]_adj_1 (BUS_ADDR_INTERNAL[1]), .n17384(n17384), 
        .\BUS_req[2] (BUS_req[2]), .\BUS_ADDR_INTERNAL[18] (BUS_ADDR_INTERNAL_adj_2610[18]), 
        .n2642(n2642), .LOGIC_CLOCK_enable_52(LOGIC_CLOCK_enable_52), .n2504(n2504), 
        .n17279(n17279), .PIC_DATA_IN_out_0(PIC_DATA_IN_out_0), .WRITE_DONE(WRITE_DONE_adj_2554), 
        .n18280(n18280), .PIC_ADDR_IN_c_1(PIC_ADDR_IN_c_1), .PIC_ADDR_IN_c_2(PIC_ADDR_IN_c_2), 
        .PIC_ADDR_IN_c_3(PIC_ADDR_IN_c_3), .PIC_ADDR_IN_c_4(PIC_ADDR_IN_c_4), 
        .PIC_ADDR_IN_c_5(PIC_ADDR_IN_c_5), .PIC_ADDR_IN_c_6(PIC_ADDR_IN_c_6), 
        .PIC_ADDR_IN_c_7(PIC_ADDR_IN_c_7), .PIC_ADDR_IN_c_8(PIC_ADDR_IN_c_8), 
        .PIC_ADDR_IN_c_9(PIC_ADDR_IN_c_9), .PIC_ADDR_IN_c_10(PIC_ADDR_IN_c_10), 
        .PIC_ADDR_IN_c_11(PIC_ADDR_IN_c_11), .PIC_ADDR_IN_c_12(PIC_ADDR_IN_c_12), 
        .PIC_ADDR_IN_c_13(PIC_ADDR_IN_c_13), .PIC_ADDR_IN_c_14(PIC_ADDR_IN_c_14), 
        .PIC_ADDR_IN_c_15(PIC_ADDR_IN_c_15), .PIC_ADDR_IN_c_16(PIC_ADDR_IN_c_16), 
        .PIC_ADDR_IN_c_17(PIC_ADDR_IN_c_17), .PIC_ADDR_IN_c_18(PIC_ADDR_IN_c_18), 
        .n14(n14), .n17434(n17434), .BUS_DIRECTION_INTERNAL(BUS_DIRECTION_INTERNAL), 
        .n18260(n18260), .n16456(n16456), .n17276(n17276), .LOGIC_CLOCK_N_57_enable_3(LOGIC_CLOCK_N_57_enable_3), 
        .n17457(n17457), .n17278(n17278), .n15571(n15571), .PIC_OE_c(PIC_OE_c), 
        .n15469(n15469), .PIC_READY_c(PIC_READY_c), .SpriteRead_yInSprite({SpriteRead_yInSprite}), 
        .\currSprite_size[6] (currSprite_size[6]), .\currSprite_size[4] (currSprite_size[4]), 
        .\currSprite_size[2] (currSprite_size[2]), .n17394(n17394), .\Sprite_readAddr_13__N_752[0] (Sprite_readAddr_13__N_752[0]), 
        .\Sprite_readAddr_13__N_752[2] (Sprite_readAddr_13__N_752[2]), .\Sprite_readAddr_13__N_752[3] (Sprite_readAddr_13__N_752[3]), 
        .\Sprite_readAddr_13__N_752[4] (Sprite_readAddr_13__N_752[4]), .\Sprite_readAddr_13__N_752[6] (Sprite_readAddr_13__N_752[6]), 
        .\Sprite_readAddr_13__N_752[5] (Sprite_readAddr_13__N_752[5]), .\Sprite_readAddr_13__N_752[8] (Sprite_readAddr_13__N_752[8]), 
        .\Sprite_readAddr_13__N_752[7] (Sprite_readAddr_13__N_752[7]), .\Sprite_readAddr_13__N_752[10] (Sprite_readAddr_13__N_752[10]), 
        .\Sprite_readAddr_13__N_752[9] (Sprite_readAddr_13__N_752[9]), .\Sprite_readAddr_13__N_752[12] (Sprite_readAddr_13__N_752[12]), 
        .\Sprite_readAddr_13__N_752[11] (Sprite_readAddr_13__N_752[11]), .\Sprite_readAddr_13__N_752[13] (Sprite_readAddr_13__N_752[13]), 
        .\currSprite_size[1] (currSprite_size[1]), .\Sprite_readAddr_13__N_752[1] (Sprite_readAddr_13__N_752[1]), 
        .\currSprite_size[3] (currSprite_size[3]), .\currSprite_size[5] (currSprite_size[5]), 
        .\currSprite_size[7] (currSprite_size[7]), .\BUS_data[1] (BUS_data[1]), 
        .\BUS_data[2] (BUS_data[2]), .\BUS_data[3] (BUS_data[3]), .\BUS_ADDR_INTERNAL[2] (BUS_ADDR_INTERNAL_adj_2610[2]), 
        .\BUS_ADDR_INTERNAL[3] (BUS_ADDR_INTERNAL_adj_2610[3]), .\BUS_ADDR_INTERNAL[4] (BUS_ADDR_INTERNAL_adj_2610[4]), 
        .\BUS_ADDR_INTERNAL[5] (BUS_ADDR_INTERNAL_adj_2610[5]), .\BUS_ADDR_INTERNAL[6] (BUS_ADDR_INTERNAL_adj_2610[6]), 
        .\BUS_ADDR_INTERNAL[7] (BUS_ADDR_INTERNAL_adj_2610[7]), .\BUS_ADDR_INTERNAL[13] (BUS_ADDR_INTERNAL_adj_2610[13]), 
        .\BUS_ADDR_INTERNAL[14] (BUS_ADDR_INTERNAL_adj_2610[14]), .\BUS_ADDR_INTERNAL[15] (BUS_ADDR_INTERNAL_adj_2610[15]), 
        .\BUS_ADDR_INTERNAL[16] (BUS_ADDR_INTERNAL_adj_2610[16]), .\BUS_ADDR_INTERNAL[17] (BUS_ADDR_INTERNAL_adj_2610[17]), 
        .\BUS_data[4] (BUS_data[4]), .\BUS_data[5] (BUS_data[5]), .\BUS_data[6] (BUS_data[6]), 
        .\BUS_data[7] (BUS_data[7]), .\writeData[4] (writeData[4]), .\writeData[5] (writeData[5]), 
        .\writeData[6] (writeData[6]), .\writeData[7] (writeData[7]), .PIC_DATA_IN_out_2(PIC_DATA_IN_out_2), 
        .PIC_DATA_IN_out_1(PIC_DATA_IN_out_1), .PIC_DATA_IN_out_4(PIC_DATA_IN_out_4), 
        .PIC_DATA_IN_out_3(PIC_DATA_IN_out_3), .PIC_DATA_IN_out_6(PIC_DATA_IN_out_6), 
        .PIC_DATA_IN_out_5(PIC_DATA_IN_out_5), .n18264(n18264), .lastAddress_31__N_1310(lastAddress_31__N_1310), 
        .n18271(n18271), .n18277(n18277), .n18266(n18266), .n18262(n18262), 
        .n18274(n18274), .n18265(n18265), .n18276(n18276), .n17409(n17409), 
        .n18275(n18275), .n17423(n17423), .n18263(n18263), .n18261(n18261), 
        .n17275(n17275), .\BUS_DATA_INTERNAL[1] (BUS_DATA_INTERNAL_adj_2609[1]), 
        .\BUS_DATA_INTERNAL[2] (BUS_DATA_INTERNAL_adj_2609[2]), .\BUS_DATA_INTERNAL[3] (BUS_DATA_INTERNAL_adj_2609[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(218[21:36])
    LUT4 m1_lut (.Z(n18280)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i12108_3_lut_4_lut (.A(n17374), .B(n17458), .C(n4266), .D(n4250), 
         .Z(n15770)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(108[14:81])
    defparam i12108_3_lut_4_lut.init = 16'hf4b0;
    
endmodule
//
// Verilog Description of module SRAM
//

module SRAM (LOGIC_CLOCK, lastAddress_31__N_1323, n66, lastAddress_31__N_1386, 
            lastAddress_31__N_1324, lastAddress_31__N_1389, lastAddress_31__N_1377, 
            lastAddress_31__N_1310, lastAddress_31__N_1325, lastAddress_31__N_1392, 
            lastAddress_31__N_1326, lastAddress_31__N_1395, lastAddress_31__N_1327, 
            lastAddress_31__N_1398, BUS_DATA_INTERNAL, n17336, SRAM_DATA_out_0, 
            lastAddress_31__N_1328, lastAddress_31__N_1401, lastAddress_31__N_1329, 
            lastAddress, lastAddress_31__N_1410, n56, SRAM_ADDR_c_0, 
            n17343, lastAddress_31__N_1332, n39, lastAddress_31__N_1339, 
            lastAddress_31__N_1431, n18280, lastAddress_31__N_1380, n46, 
            lastAddress_31__N_1416, n58, n45, lastAddress_31__N_1434, 
            n64, \BUS_ADDR_INTERNAL[18]_derived_1 , lastAddress_31__N_1334, 
            BUS_DONE_INTERNAL, SRAM_WE_N_1254, \BUS_addr[10] , lastAddress_31__N_1404, 
            \lastAddress[7] , lastAddress_31__N_1413, n57, lastAddress_31__N_1419, 
            n59, n40, \lastAddress[5] , \lastAddress[24] , SRAM_OE_c, 
            SRAM_WE_c, lastAddress_31__N_1335, n41, n18260, n42, lastAddress_31__N_1422, 
            n60, n43, lastAddress_31__N_1340, lastAddress_31__N_1336, 
            n4, \BUS_data[9] , \lastAddress[23] , n4_adj_22, \BUS_data[10] , 
            n4_adj_23, \BUS_data[11] , n4_adj_24, \BUS_data[12] , n4_adj_25, 
            \BUS_data[13] , n4_adj_26, \BUS_data[14] , lastAddress_31__N_1425, 
            n61, n4_adj_27, \BUS_data[15] , \lastAddress[22] , n4_adj_28, 
            \BUS_data[4] , \lastAddress[4] , n4_adj_29, \BUS_data[5] , 
            n4_adj_30, \BUS_data[6] , lastAddress_31__N_1337, n4_adj_31, 
            \BUS_data[7] , lastAddress_31__N_1383, lastAddress_31__N_1428, 
            n62, \lastAddress[30] , n33, n35, \lastAddress[21] , lastAddress_31__N_1338, 
            \BUS_DATA_INTERNAL[1] , SRAM_DATA_out_1, \BUS_DATA_INTERNAL[2] , 
            SRAM_DATA_out_2, \BUS_DATA_INTERNAL[3] , SRAM_DATA_out_3, 
            SRAM_DATA_out_4, SRAM_DATA_out_5, SRAM_DATA_out_6, SRAM_DATA_out_7, 
            \BUS_DATA_INTERNAL[8] , SRAM_DATA_out_8, SRAM_DATA_out_9, 
            SRAM_DATA_out_10, SRAM_DATA_out_11, SRAM_DATA_out_12, SRAM_DATA_out_13, 
            SRAM_DATA_out_14, SRAM_DATA_out_15, lastAddress_31__N_1333, 
            n36, \lastAddress[3] , \lastAddress[20] , SRAM_ADDR_c_1, 
            n17342, SRAM_ADDR_c_2, n17339, SRAM_ADDR_c_3, n17333, 
            SRAM_ADDR_c_4, n17332, SRAM_ADDR_c_5, n17331, SRAM_ADDR_c_6, 
            n17321, SRAM_ADDR_c_7, n17334, SRAM_ADDR_c_8, n17337, 
            SRAM_ADDR_c_9, n17325, SRAM_ADDR_c_10, SRAM_ADDR_c_11, \BUS_addr[11] , 
            SRAM_ADDR_c_12, n17335, SRAM_ADDR_c_13, n17338, SRAM_ADDR_c_14, 
            n17322, SRAM_ADDR_c_15, n17320, SRAM_ADDR_c_16, n17323, 
            SRAM_ADDR_c_17, n17340, lastAddress_31__N_1331, lastAddress_31__N_1407, 
            lastAddress_31__N_1330, \lastAddress[2] , \lastAddress[31] , 
            n63, \lastAddress[17] , \lastAddress[29] , \lastAddress[13] , 
            \lastAddress[12] , GND_net, \lastAddress[16] , \lastAddress[15] , 
            \lastAddress[14] , \lastAddress[28] , \lastAddress[27] , \lastAddress[26] , 
            \lastAddress[1] , n55, \lastAddress[9] , n17287, n7, n9, 
            n6250, \lastAddress[8] );
    input LOGIC_CLOCK;
    input lastAddress_31__N_1323;
    input [31:0]n66;
    input lastAddress_31__N_1386;
    input lastAddress_31__N_1324;
    input lastAddress_31__N_1389;
    input lastAddress_31__N_1377;
    input lastAddress_31__N_1310;
    input lastAddress_31__N_1325;
    input lastAddress_31__N_1392;
    input lastAddress_31__N_1326;
    input lastAddress_31__N_1395;
    input lastAddress_31__N_1327;
    input lastAddress_31__N_1398;
    output [15:0]BUS_DATA_INTERNAL;
    input n17336;
    input SRAM_DATA_out_0;
    input lastAddress_31__N_1328;
    input lastAddress_31__N_1401;
    input lastAddress_31__N_1329;
    output [31:0]lastAddress;
    input lastAddress_31__N_1410;
    input n56;
    output SRAM_ADDR_c_0;
    input n17343;
    input lastAddress_31__N_1332;
    input n39;
    input lastAddress_31__N_1339;
    input lastAddress_31__N_1431;
    input n18280;
    input lastAddress_31__N_1380;
    input n46;
    input lastAddress_31__N_1416;
    input n58;
    input n45;
    input lastAddress_31__N_1434;
    input n64;
    input \BUS_ADDR_INTERNAL[18]_derived_1 ;
    input lastAddress_31__N_1334;
    output BUS_DONE_INTERNAL;
    output SRAM_WE_N_1254;
    input \BUS_addr[10] ;
    input lastAddress_31__N_1404;
    output \lastAddress[7] ;
    input lastAddress_31__N_1413;
    input n57;
    input lastAddress_31__N_1419;
    input n59;
    input n40;
    output \lastAddress[5] ;
    output \lastAddress[24] ;
    output SRAM_OE_c;
    output SRAM_WE_c;
    input lastAddress_31__N_1335;
    input n41;
    input n18260;
    input n42;
    input lastAddress_31__N_1422;
    input n60;
    input n43;
    input lastAddress_31__N_1340;
    input lastAddress_31__N_1336;
    input n4;
    output \BUS_data[9] ;
    output \lastAddress[23] ;
    input n4_adj_22;
    output \BUS_data[10] ;
    input n4_adj_23;
    output \BUS_data[11] ;
    input n4_adj_24;
    output \BUS_data[12] ;
    input n4_adj_25;
    output \BUS_data[13] ;
    input n4_adj_26;
    output \BUS_data[14] ;
    input lastAddress_31__N_1425;
    input n61;
    input n4_adj_27;
    output \BUS_data[15] ;
    output \lastAddress[22] ;
    input n4_adj_28;
    output \BUS_data[4] ;
    output \lastAddress[4] ;
    input n4_adj_29;
    output \BUS_data[5] ;
    input n4_adj_30;
    output \BUS_data[6] ;
    input lastAddress_31__N_1337;
    input n4_adj_31;
    output \BUS_data[7] ;
    input lastAddress_31__N_1383;
    input lastAddress_31__N_1428;
    input n62;
    output \lastAddress[30] ;
    input n33;
    input n35;
    output \lastAddress[21] ;
    input lastAddress_31__N_1338;
    output \BUS_DATA_INTERNAL[1] ;
    input SRAM_DATA_out_1;
    output \BUS_DATA_INTERNAL[2] ;
    input SRAM_DATA_out_2;
    output \BUS_DATA_INTERNAL[3] ;
    input SRAM_DATA_out_3;
    input SRAM_DATA_out_4;
    input SRAM_DATA_out_5;
    input SRAM_DATA_out_6;
    input SRAM_DATA_out_7;
    output \BUS_DATA_INTERNAL[8] ;
    input SRAM_DATA_out_8;
    input SRAM_DATA_out_9;
    input SRAM_DATA_out_10;
    input SRAM_DATA_out_11;
    input SRAM_DATA_out_12;
    input SRAM_DATA_out_13;
    input SRAM_DATA_out_14;
    input SRAM_DATA_out_15;
    input lastAddress_31__N_1333;
    input n36;
    output \lastAddress[3] ;
    output \lastAddress[20] ;
    output SRAM_ADDR_c_1;
    input n17342;
    output SRAM_ADDR_c_2;
    input n17339;
    output SRAM_ADDR_c_3;
    input n17333;
    output SRAM_ADDR_c_4;
    input n17332;
    output SRAM_ADDR_c_5;
    input n17331;
    output SRAM_ADDR_c_6;
    input n17321;
    output SRAM_ADDR_c_7;
    input n17334;
    output SRAM_ADDR_c_8;
    input n17337;
    output SRAM_ADDR_c_9;
    input n17325;
    output SRAM_ADDR_c_10;
    output SRAM_ADDR_c_11;
    input \BUS_addr[11] ;
    output SRAM_ADDR_c_12;
    input n17335;
    output SRAM_ADDR_c_13;
    input n17338;
    output SRAM_ADDR_c_14;
    input n17322;
    output SRAM_ADDR_c_15;
    input n17320;
    output SRAM_ADDR_c_16;
    input n17323;
    output SRAM_ADDR_c_17;
    input n17340;
    input lastAddress_31__N_1331;
    input lastAddress_31__N_1407;
    input lastAddress_31__N_1330;
    output \lastAddress[2] ;
    output \lastAddress[31] ;
    input n63;
    output \lastAddress[17] ;
    output \lastAddress[29] ;
    output \lastAddress[13] ;
    output \lastAddress[12] ;
    input GND_net;
    output \lastAddress[16] ;
    output \lastAddress[15] ;
    output \lastAddress[14] ;
    output \lastAddress[28] ;
    output \lastAddress[27] ;
    output \lastAddress[26] ;
    output \lastAddress[1] ;
    input n55;
    output \lastAddress[9] ;
    input n17287;
    input n7;
    input n9;
    output n6250;
    output \lastAddress[8] ;
    
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    
    wire n7123, n7120, n7119, n7116, n7132, n7131, n7138, n7159, 
        n7156, n7115, n7112, n7111, n7108, n7107, n7104, SRAM_OE_N_1511, 
        n7103, n7100;
    wire [31:0]n66_c;
    
    wire n7099, n7153, n7152, n7130, n7088, LOGIC_CLOCK_enable_213, 
        n7087;
    wire [7:0]state;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(34[8:13])
    wire [7:0]state_7__N_1453;
    
    wire n7058, n7128, n6, n49_adj_2509, n51_adj_2510, n7127, n7126, 
        n7080, n7135, n7056, n7079, n3816, n7078, n7134, n7055, 
        n7054, n17346;
    wire [31:0]lastAddress_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(29[8:19])
    
    wire n7096, n7095, n7094, n17469, n11, n7084, n7083, n7082, 
        n7076, n7150, n7075, n7074, n7149, n5990, LOGIC_CLOCK_enable_46, 
        LOGIC_CLOCK_enable_47, SRAM_WE_N_1245, n7147, n17440, n17395, 
        n15334, n17356, n17005, n7144, n7072, n7141, n7071;
    wire [15:0]BUS_DATA_INTERNAL_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(30[8:25])
    
    wire n7146, n7068, n7143, n7070, n7067, n7124, n7064, n7168, 
        n17006, n7165, n17455, n7140, n7063, n22, n7162, n7066, 
        n7137, n7062, n7086, n7090, n7098, n7102, n7106, n7110, 
        n7114, n7118, n7122, n7155, n7158, n7161, n7164, n7167, 
        n7060, n13657, n13658, n13662, n13656, n13661, n13660, 
        n13659, n7092, n7091, n7059, n17432, n17345, n4_adj_2521, 
        n23, n19, n20, n20_adj_2522, n17319, n17007, n17282;
    wire [7:0]state_7__N_1461;
    
    FD1S3BX lastAddress_i0_i17_3771_3772_set (.D(n66[17]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1323), .Q(n7123)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i17_3771_3772_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i16_3767_3768_reset (.D(n66[16]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1386), .Q(n7120)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i16_3767_3768_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i16_3767_3768_set (.D(n66[16]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1324), .Q(n7119)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i16_3767_3768_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i15_3763_3764_reset (.D(n66[15]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1389), .Q(n7116)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i15_3763_3764_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i30_3779_3780_reset (.D(n66[30]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7132)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i30_3779_3780_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i30_3779_3780_set (.D(n66[30]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7131)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i30_3779_3780_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i20_3785_3786_reset (.D(n66[20]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7138)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i20_3785_3786_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i27_3806_3807_reset (.D(n66[27]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7159)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i27_3806_3807_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i26_3803_3804_reset (.D(n66[26]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7156)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i26_3803_3804_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i15_3763_3764_set (.D(n66[15]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1325), .Q(n7115)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i15_3763_3764_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i14_3759_3760_reset (.D(n66[14]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1392), .Q(n7112)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i14_3759_3760_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i14_3759_3760_set (.D(n66[14]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1326), .Q(n7111)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i14_3759_3760_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i13_3755_3756_reset (.D(n66[13]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1395), .Q(n7108)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i13_3755_3756_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i13_3755_3756_set (.D(n66[13]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1327), .Q(n7107)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i13_3755_3756_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i12_3751_3752_reset (.D(n66[12]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1398), .Q(n7104)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i12_3751_3752_reset.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i0 (.D(SRAM_DATA_out_0), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i0.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i12_3751_3752_set (.D(n66[12]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1328), .Q(n7103)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i12_3751_3752_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i11_3747_3748_reset (.D(n66_c[11]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1401), .Q(n7100)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i11_3747_3748_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i11_3747_3748_set (.D(n66_c[11]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1329), .Q(n7099)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i11_3747_3748_set.GSR = "DISABLED";
    LUT4 i3802_3_lut (.A(n7153), .B(n7152), .C(n7130), .Z(lastAddress[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3802_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i8_3735_3736_reset (.D(n56), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1410), .Q(n7088)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i8_3735_3736_reset.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i1 (.D(n17343), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i1.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i8_3735_3736_set (.D(n56), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1332), .Q(n7087)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i8_3735_3736_set.GSR = "DISABLED";
    FD1S3DX state_i0 (.D(state_7__N_1453[0]), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam state_i0.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i25_3800_3801_reset (.D(n39), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7153)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i25_3800_3801_reset.GSR = "DISABLED";
    FD1S1D i3706 (.D(n18280), .CK(lastAddress_31__N_1339), .CD(lastAddress_31__N_1431), 
           .Q(n7058));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3706.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i18_3775_3776_reset (.D(n46), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1380), .Q(n7128)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i18_3775_3776_reset.GSR = "DISABLED";
    PFUMX i55 (.BLUT(n6), .ALUT(n49_adj_2509), .C0(state[4]), .Z(n51_adj_2510));
    LUT4 i3777_3_lut (.A(n7128), .B(n7127), .C(n7126), .Z(lastAddress[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3777_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i6_3727_3728_reset (.D(n58), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1416), .Q(n7080)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i6_3727_3728_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i19_3782_3783_reset (.D(n45), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7135)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i19_3782_3783_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i0_3703_3704_reset (.D(n64), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1434), .Q(n7056)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i0_3703_3704_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i18_3775_3776_set (.D(n46), .CK(LOGIC_CLOCK), 
            .PD(\BUS_ADDR_INTERNAL[18]_derived_1 ), .Q(n7127)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i18_3775_3776_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i6_3727_3728_set (.D(n58), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1334), .Q(n7079)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i6_3727_3728_set.GSR = "DISABLED";
    FD1S3DX BUS_DONE_INTERNAL_128 (.D(n3816), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(BUS_DONE_INTERNAL)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DONE_INTERNAL_128.GSR = "DISABLED";
    LUT4 i3729_3_lut (.A(n7080), .B(n7079), .C(n7078), .Z(lastAddress[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3729_3_lut.init = 16'hcaca;
    LUT4 i3784_3_lut (.A(n7135), .B(n7134), .C(n7130), .Z(lastAddress[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3784_3_lut.init = 16'hcaca;
    LUT4 i3705_3_lut (.A(n7056), .B(n7055), .C(n7054), .Z(lastAddress[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3705_3_lut.init = 16'hcaca;
    LUT4 i6600_3_lut (.A(BUS_DONE_INTERNAL), .B(SRAM_WE_N_1254), .C(n17346), 
         .Z(n3816)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i6600_3_lut.init = 16'h8c8c;
    LUT4 lastAddress_i1_i11_3_lut (.A(lastAddress_c[10]), .B(\BUS_addr[10] ), 
         .C(SRAM_WE_N_1254), .Z(n66_c[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i1_i11_3_lut.init = 16'hacac;
    LUT4 i3745_3_lut (.A(n7096), .B(n7095), .C(n7094), .Z(lastAddress_c[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3745_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(n17469), .C(state[5]), .D(state[4]), 
         .Z(n11)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_3_lut_4_lut.init = 16'hf8f0;
    FD1S3DX lastAddress_i0_i10_3743_3744_reset (.D(n66_c[10]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1404), .Q(n7096)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i10_3743_3744_reset.GSR = "DISABLED";
    LUT4 i3733_3_lut (.A(n7084), .B(n7083), .C(n7082), .Z(\lastAddress[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3733_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i7_3731_3732_reset (.D(n57), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1413), .Q(n7084)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i7_3731_3732_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i5_3723_3724_reset (.D(n59), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1419), .Q(n7076)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i5_3723_3724_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i24_3797_3798_reset (.D(n40), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7150)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i24_3797_3798_reset.GSR = "DISABLED";
    LUT4 i3725_3_lut (.A(n7076), .B(n7075), .C(n7074), .Z(\lastAddress[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3725_3_lut.init = 16'hcaca;
    LUT4 i3799_3_lut (.A(n7150), .B(n7149), .C(n7130), .Z(\lastAddress[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3799_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(state[5]), .B(state[1]), .C(state[2]), .D(state[3]), 
         .Z(n5990)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hbfff;
    FD1P3BX SRAM_OE_INT_230 (.D(SRAM_OE_N_1511), .SP(LOGIC_CLOCK_enable_46), 
            .CK(LOGIC_CLOCK), .PD(n17336), .Q(SRAM_OE_c)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_OE_INT_230.GSR = "DISABLED";
    FD1P3BX SRAM_WE_INT_229 (.D(SRAM_WE_N_1245), .SP(LOGIC_CLOCK_enable_47), 
            .CK(LOGIC_CLOCK), .PD(n17336), .Q(SRAM_WE_c)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_WE_INT_229.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i5_3723_3724_set (.D(n59), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1335), .Q(n7075)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i5_3723_3724_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i23_3794_3795_reset (.D(n41), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7147)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i23_3794_3795_reset.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_432 (.A(state[1]), .B(state[2]), .Z(n17440)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_2_lut_rep_432.init = 16'heeee;
    LUT4 i1_2_lut_rep_387_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n17395)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_2_lut_rep_387_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n18260), 
         .D(state[0]), .Z(n15334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_348_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[0]), .Z(n17356)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_2_lut_rep_348_3_lut_4_lut.init = 16'hfffe;
    LUT4 state_7__N_1469_0__bdd_4_lut_13265 (.A(state[0]), .B(state[3]), 
         .C(state[2]), .D(state[1]), .Z(n17005)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam state_7__N_1469_0__bdd_4_lut_13265.init = 16'h4000;
    FD1S3DX lastAddress_i0_i22_3791_3792_reset (.D(n42), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7144)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i22_3791_3792_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i4_3719_3720_reset (.D(n60), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1422), .Q(n7072)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i4_3719_3720_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i21_3788_3789_reset (.D(n43), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7141)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i21_3788_3789_reset.GSR = "DISABLED";
    FD1S1D i3702 (.D(n18280), .CK(lastAddress_31__N_1340), .CD(lastAddress_31__N_1434), 
           .Q(n7054));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3702.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i4_3719_3720_set (.D(n60), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1336), .Q(n7071)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i4_3719_3720_set.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_adj_657 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4), .D(BUS_DATA_INTERNAL_c[9]), .Z(\BUS_data[9] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_657.init = 16'hf4f0;
    LUT4 i3796_3_lut (.A(n7147), .B(n7146), .C(n7130), .Z(\lastAddress[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3796_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_adj_658 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_22), .D(BUS_DATA_INTERNAL_c[10]), .Z(\BUS_data[10] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_658.init = 16'hf4f0;
    LUT4 i2_3_lut_4_lut_adj_659 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_23), .D(BUS_DATA_INTERNAL_c[11]), .Z(\BUS_data[11] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_659.init = 16'hf4f0;
    LUT4 i2_3_lut_4_lut_adj_660 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_24), .D(BUS_DATA_INTERNAL_c[12]), .Z(\BUS_data[12] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_660.init = 16'hf4f0;
    LUT4 i2_3_lut_4_lut_adj_661 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_25), .D(BUS_DATA_INTERNAL_c[13]), .Z(\BUS_data[13] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_661.init = 16'hf4f0;
    LUT4 i2_3_lut_4_lut_adj_662 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_26), .D(BUS_DATA_INTERNAL_c[14]), .Z(\BUS_data[14] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_662.init = 16'hf4f0;
    FD1S3DX lastAddress_i0_i3_3715_3716_reset (.D(n61), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1425), .Q(n7068)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i3_3715_3716_reset.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_adj_663 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_27), .D(BUS_DATA_INTERNAL_c[15]), .Z(\BUS_data[15] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_663.init = 16'hf4f0;
    LUT4 i3793_3_lut (.A(n7144), .B(n7143), .C(n7130), .Z(\lastAddress[22] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3793_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_adj_664 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_28), .D(BUS_DATA_INTERNAL_c[4]), .Z(\BUS_data[4] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_664.init = 16'hf4f0;
    LUT4 i3721_3_lut (.A(n7072), .B(n7071), .C(n7070), .Z(\lastAddress[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3721_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_adj_665 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_29), .D(BUS_DATA_INTERNAL_c[5]), .Z(\BUS_data[5] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_665.init = 16'hf4f0;
    LUT4 i2_3_lut_4_lut_adj_666 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_30), .D(BUS_DATA_INTERNAL_c[6]), .Z(\BUS_data[6] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_666.init = 16'hf4f0;
    FD1S3BX lastAddress_i0_i3_3715_3716_set (.D(n61), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1337), .Q(n7067)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i3_3715_3716_set.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_adj_667 (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n18260), 
         .C(n4_adj_31), .D(BUS_DATA_INTERNAL_c[7]), .Z(\BUS_data[7] )) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(45[41:88])
    defparam i2_3_lut_4_lut_adj_667.init = 16'hf4f0;
    FD1S3DX lastAddress_i0_i17_3771_3772_reset (.D(n66[17]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1383), .Q(n7124)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i17_3771_3772_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i2_3711_3712_reset (.D(n62), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1428), .Q(n7064)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i2_3711_3712_reset.GSR = "DISABLED";
    LUT4 i3781_3_lut (.A(n7132), .B(n7131), .C(n7130), .Z(\lastAddress[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3781_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i31_3815_3816_reset (.D(n33), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7168)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i31_3815_3816_reset.GSR = "DISABLED";
    LUT4 state_7__N_1469_0__bdd_4_lut (.A(n18260), .B(state[3]), .C(state[2]), 
         .D(state[1]), .Z(n17006)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam state_7__N_1469_0__bdd_4_lut.init = 16'h0002;
    FD1S3BX lastAddress_i0_i0_3703_3704_set (.D(n64), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1340), .Q(n7055)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i0_3703_3704_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i29_3812_3813_reset (.D(n35), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7165)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i29_3812_3813_reset.GSR = "DISABLED";
    LUT4 i2_3_lut_rep_447 (.A(state[4]), .B(state[5]), .C(state[0]), .Z(n17455)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i2_3_lut_rep_447.init = 16'hfefe;
    LUT4 i3790_3_lut (.A(n7141), .B(n7140), .C(n7130), .Z(\lastAddress[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3790_3_lut.init = 16'hcaca;
    FD1S3BX lastAddress_i0_i2_3711_3712_set (.D(n62), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1338), .Q(n7063)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i2_3711_3712_set.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_3_lut (.A(state[0]), .B(state[1]), .C(state[5]), 
         .Z(n22)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_2_lut_3_lut_3_lut.init = 16'hf7f7;
    FD1P3DX BUS_DATA_INTERNAL_i0_i1 (.D(SRAM_DATA_out_1), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(\BUS_DATA_INTERNAL[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i1.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i2 (.D(SRAM_DATA_out_2), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(\BUS_DATA_INTERNAL[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i2.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i3 (.D(SRAM_DATA_out_3), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(\BUS_DATA_INTERNAL[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i3.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i4 (.D(SRAM_DATA_out_4), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i4.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i5 (.D(SRAM_DATA_out_5), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i5.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i6 (.D(SRAM_DATA_out_6), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i6.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i7 (.D(SRAM_DATA_out_7), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i7.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i8 (.D(SRAM_DATA_out_8), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(\BUS_DATA_INTERNAL[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i8.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i9 (.D(SRAM_DATA_out_9), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i9.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i10 (.D(SRAM_DATA_out_10), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i10.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i11 (.D(SRAM_DATA_out_11), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i11.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i12 (.D(SRAM_DATA_out_12), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i12.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i13 (.D(SRAM_DATA_out_13), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i13.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i14 (.D(SRAM_DATA_out_14), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i14.GSR = "DISABLED";
    FD1P3DX BUS_DATA_INTERNAL_i0_i15 (.D(SRAM_DATA_out_15), .SP(SRAM_OE_N_1511), 
            .CK(LOGIC_CLOCK), .CD(n17336), .Q(BUS_DATA_INTERNAL_c[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam BUS_DATA_INTERNAL_i0_i15.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i7_3731_3732_set (.D(n57), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1333), .Q(n7083)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i7_3731_3732_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i28_3809_3810_reset (.D(n36), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1377), .Q(n7162)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i28_3809_3810_reset.GSR = "DISABLED";
    LUT4 i3717_3_lut (.A(n7068), .B(n7067), .C(n7066), .Z(\lastAddress[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3717_3_lut.init = 16'hcaca;
    LUT4 i3787_3_lut (.A(n7138), .B(n7137), .C(n7130), .Z(\lastAddress[20] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3787_3_lut.init = 16'hcaca;
    FD1P3AX SRAM_ADDR_i0_i2 (.D(n17342), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i2.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i3 (.D(n17339), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i3.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i4 (.D(n17333), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i4.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i5 (.D(n17332), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i5.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i6 (.D(n17331), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i6.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i7 (.D(n17321), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i7.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i8 (.D(n17334), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i8.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i9 (.D(n17337), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i9.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i10 (.D(n17325), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_9)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i10.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i11 (.D(\BUS_addr[10] ), .SP(LOGIC_CLOCK_enable_213), 
            .CK(LOGIC_CLOCK), .Q(SRAM_ADDR_c_10)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i11.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i12 (.D(\BUS_addr[11] ), .SP(LOGIC_CLOCK_enable_213), 
            .CK(LOGIC_CLOCK), .Q(SRAM_ADDR_c_11)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i12.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i13 (.D(n17335), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_12)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i13.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i14 (.D(n17338), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_13)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i14.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i15 (.D(n17322), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_14)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i15.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i16 (.D(n17320), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_15)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i16.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i17 (.D(n17323), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_16)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i17.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i18 (.D(n17340), .SP(LOGIC_CLOCK_enable_213), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_17)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam SRAM_ADDR_i0_i18.GSR = "DISABLED";
    FD1S3DX state_i1 (.D(state_7__N_1453[1]), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam state_i1.GSR = "DISABLED";
    FD1S3DX state_i2 (.D(state_7__N_1453[2]), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam state_i2.GSR = "DISABLED";
    FD1S3DX state_i3 (.D(state_7__N_1453[3]), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam state_i3.GSR = "DISABLED";
    FD1S3DX state_i4 (.D(state_7__N_1453[4]), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam state_i4.GSR = "DISABLED";
    FD1S3DX state_i5 (.D(state_7__N_1453[5]), .CK(LOGIC_CLOCK), .CD(n17336), 
            .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam state_i5.GSR = "DISABLED";
    FD1S1D i3710 (.D(n18280), .CK(lastAddress_31__N_1338), .CD(lastAddress_31__N_1428), 
           .Q(n7062));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3710.GSR = "DISABLED";
    FD1S1D i3714 (.D(n18280), .CK(lastAddress_31__N_1337), .CD(lastAddress_31__N_1425), 
           .Q(n7066));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3714.GSR = "DISABLED";
    FD1S1D i3718 (.D(n18280), .CK(lastAddress_31__N_1336), .CD(lastAddress_31__N_1422), 
           .Q(n7070));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3718.GSR = "DISABLED";
    FD1S1D i3722 (.D(n18280), .CK(lastAddress_31__N_1335), .CD(lastAddress_31__N_1419), 
           .Q(n7074));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3722.GSR = "DISABLED";
    FD1S1D i3726 (.D(n18280), .CK(lastAddress_31__N_1334), .CD(lastAddress_31__N_1416), 
           .Q(n7078));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3726.GSR = "DISABLED";
    FD1S1D i3730 (.D(n18280), .CK(lastAddress_31__N_1333), .CD(lastAddress_31__N_1413), 
           .Q(n7082));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3730.GSR = "DISABLED";
    FD1S1D i3734 (.D(n18280), .CK(lastAddress_31__N_1332), .CD(lastAddress_31__N_1410), 
           .Q(n7086));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3734.GSR = "DISABLED";
    FD1S1D i3738 (.D(n18280), .CK(lastAddress_31__N_1331), .CD(lastAddress_31__N_1407), 
           .Q(n7090));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3738.GSR = "DISABLED";
    FD1S1D i3742 (.D(n18280), .CK(lastAddress_31__N_1330), .CD(lastAddress_31__N_1404), 
           .Q(n7094));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3742.GSR = "DISABLED";
    FD1S1D i3746 (.D(n18280), .CK(lastAddress_31__N_1329), .CD(lastAddress_31__N_1401), 
           .Q(n7098));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3746.GSR = "DISABLED";
    FD1S1D i3750 (.D(n18280), .CK(lastAddress_31__N_1328), .CD(lastAddress_31__N_1398), 
           .Q(n7102));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3750.GSR = "DISABLED";
    FD1S1D i3754 (.D(n18280), .CK(lastAddress_31__N_1327), .CD(lastAddress_31__N_1395), 
           .Q(n7106));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3754.GSR = "DISABLED";
    FD1S1D i3758 (.D(n18280), .CK(lastAddress_31__N_1326), .CD(lastAddress_31__N_1392), 
           .Q(n7110));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3758.GSR = "DISABLED";
    FD1S1D i3762 (.D(n18280), .CK(lastAddress_31__N_1325), .CD(lastAddress_31__N_1389), 
           .Q(n7114));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3762.GSR = "DISABLED";
    FD1S1D i3766 (.D(n18280), .CK(lastAddress_31__N_1324), .CD(lastAddress_31__N_1386), 
           .Q(n7118));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3766.GSR = "DISABLED";
    FD1S1D i3770 (.D(n18280), .CK(lastAddress_31__N_1323), .CD(lastAddress_31__N_1383), 
           .Q(n7122));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3770.GSR = "DISABLED";
    FD1S1D i3774 (.D(n18280), .CK(\BUS_ADDR_INTERNAL[18]_derived_1 ), .CD(lastAddress_31__N_1380), 
           .Q(n7126));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3774.GSR = "DISABLED";
    FD1S1D i3778 (.D(n18280), .CK(lastAddress_31__N_1310), .CD(lastAddress_31__N_1377), 
           .Q(n7130));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3778.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i20_3785_3786_set (.D(n66[20]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7137)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i20_3785_3786_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i21_3788_3789_set (.D(n43), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7140)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i21_3788_3789_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i22_3791_3792_set (.D(n42), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7143)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i22_3791_3792_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i23_3794_3795_set (.D(n41), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7146)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i23_3794_3795_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i24_3797_3798_set (.D(n40), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7149)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i24_3797_3798_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i25_3800_3801_set (.D(n39), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7152)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i25_3800_3801_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i26_3803_3804_set (.D(n66[26]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7155)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i26_3803_3804_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i27_3806_3807_set (.D(n66[27]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7158)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i27_3806_3807_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i28_3809_3810_set (.D(n36), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7161)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i28_3809_3810_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i29_3812_3813_set (.D(n35), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7164)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i29_3812_3813_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i31_3815_3816_set (.D(n33), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7167)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i31_3815_3816_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i19_3782_3783_set (.D(n45), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1310), .Q(n7134)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i19_3782_3783_set.GSR = "DISABLED";
    LUT4 i3713_3_lut (.A(n7064), .B(n7063), .C(n7062), .Z(\lastAddress[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3713_3_lut.init = 16'hcaca;
    LUT4 i3817_3_lut (.A(n7168), .B(n7167), .C(n7130), .Z(\lastAddress[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3817_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i1_3707_3708_reset (.D(n63), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1431), .Q(n7060)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i1_3707_3708_reset.GSR = "DISABLED";
    LUT4 i3773_3_lut (.A(n7124), .B(n7123), .C(n7122), .Z(\lastAddress[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3773_3_lut.init = 16'hcaca;
    LUT4 i3814_3_lut (.A(n7165), .B(n7164), .C(n7130), .Z(\lastAddress[29] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3814_3_lut.init = 16'hcaca;
    CCU2D lastAddress_31__I_0_304_23 (.A0(n17338), .B0(\lastAddress[13] ), 
          .C0(n17335), .D0(\lastAddress[12] ), .A1(\BUS_addr[11] ), .B1(lastAddress_c[11]), 
          .C1(\BUS_addr[10] ), .D1(lastAddress_c[10]), .CIN(n13657), .COUT(n13658));
    defparam lastAddress_31__I_0_304_23.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_304_23.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_304_23.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_23.INJECT1_1 = "YES";
    FD1S3BX lastAddress_i0_i10_3743_3744_set (.D(n66_c[10]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1330), .Q(n7095)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i10_3743_3744_set.GSR = "DISABLED";
    CCU2D lastAddress_31__I_0_304_32 (.A0(\lastAddress[22] ), .B0(\lastAddress[21] ), 
          .C0(\lastAddress[20] ), .D0(lastAddress[19]), .A1(GND_net), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n13662), .S1(SRAM_WE_N_1254));
    defparam lastAddress_31__I_0_304_32.INIT0 = 16'h8001;
    defparam lastAddress_31__I_0_304_32.INIT1 = 16'hFFFF;
    defparam lastAddress_31__I_0_304_32.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_32.INJECT1_1 = "NO";
    CCU2D lastAddress_31__I_0_304_21 (.A0(n17340), .B0(\lastAddress[17] ), 
          .C0(n17323), .D0(\lastAddress[16] ), .A1(n17320), .B1(\lastAddress[15] ), 
          .C1(n17322), .D1(\lastAddress[14] ), .CIN(n13656), .COUT(n13657));
    defparam lastAddress_31__I_0_304_21.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_304_21.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_304_21.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_21.INJECT1_1 = "YES";
    CCU2D lastAddress_31__I_0_304_31 (.A0(\lastAddress[28] ), .B0(\lastAddress[27] ), 
          .C0(\lastAddress[26] ), .D0(lastAddress[25]), .A1(lastAddress[25]), 
          .B1(\lastAddress[24] ), .C1(\lastAddress[23] ), .D1(\lastAddress[22] ), 
          .CIN(n13661), .COUT(n13662));
    defparam lastAddress_31__I_0_304_31.INIT0 = 16'h8001;
    defparam lastAddress_31__I_0_304_31.INIT1 = 16'h8001;
    defparam lastAddress_31__I_0_304_31.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_31.INJECT1_1 = "YES";
    CCU2D lastAddress_31__I_0_304_29 (.A0(n17342), .B0(\lastAddress[1] ), 
          .C0(n17343), .D0(lastAddress[0]), .A1(lastAddress_31__N_1310), 
          .B1(\lastAddress[30] ), .C1(\lastAddress[29] ), .D1(\lastAddress[28] ), 
          .CIN(n13660), .COUT(n13661));
    defparam lastAddress_31__I_0_304_29.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_304_29.INIT1 = 16'h8001;
    defparam lastAddress_31__I_0_304_29.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_29.INJECT1_1 = "YES";
    CCU2D lastAddress_31__I_0_304_27 (.A0(n17331), .B0(\lastAddress[5] ), 
          .C0(n17332), .D0(\lastAddress[4] ), .A1(n17333), .B1(\lastAddress[3] ), 
          .C1(n17339), .D1(\lastAddress[2] ), .CIN(n13659), .COUT(n13660));
    defparam lastAddress_31__I_0_304_27.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_304_27.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_304_27.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_27.INJECT1_1 = "YES";
    FD1S3DX lastAddress_i0_i9_3739_3740_reset (.D(n55), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_1407), .Q(n7092)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i9_3739_3740_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i9_3739_3740_set (.D(n55), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1331), .Q(n7091)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i9_3739_3740_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i1_3707_3708_set (.D(n63), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_1339), .Q(n7059)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=199, LSE_RLINE=199 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i0_i1_3707_3708_set.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_461 (.A(state[2]), .B(state[1]), .Z(n17469)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_2_lut_rep_461.init = 16'h8888;
    LUT4 i1_2_lut_rep_424_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n17432)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_2_lut_rep_424_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_rep_337_4_lut_4_lut (.A(state[5]), .B(state[4]), .C(state[3]), 
         .D(n17395), .Z(n17345)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(94[10:23])
    defparam i2_3_lut_rep_337_4_lut_4_lut.init = 16'hfffd;
    LUT4 i2_4_lut_4_lut (.A(state[5]), .B(state[3]), .C(n17432), .D(n15334), 
         .Z(n6)) /* synthesis lut_function=(!(A+!(B (C)+!B !(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(94[10:23])
    defparam i2_4_lut_4_lut.init = 16'h4051;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n17395), .B(state[3]), .C(state[5]), 
         .D(state[4]), .Z(n4_adj_2521)) /* synthesis lut_function=(A (C)+!A !(B+!(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hb1b0;
    LUT4 i1_3_lut_rep_338_4_lut (.A(n17395), .B(state[3]), .C(state[5]), 
         .D(state[4]), .Z(n17346)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_3_lut_rep_338_4_lut.init = 16'heeef;
    LUT4 i3811_3_lut (.A(n7162), .B(n7161), .C(n7130), .Z(\lastAddress[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3811_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(SRAM_WE_N_1254), .B(state[3]), .C(n23), .D(n19), 
         .Z(state_7__N_1453[1])) /* synthesis lut_function=((B (C)+!B (C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_4_lut.init = 16'hf7f5;
    LUT4 i1_4_lut_adj_668 (.A(state[1]), .B(state[5]), .C(state[2]), .D(state[0]), 
         .Z(n23)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_4_lut_adj_668.init = 16'h8aaa;
    LUT4 i1_3_lut (.A(n17455), .B(state[1]), .C(state[2]), .Z(n19)) /* synthesis lut_function=(A (B)+!A (B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_3_lut.init = 16'hcdcd;
    LUT4 i2_4_lut (.A(state[2]), .B(n20), .C(n22), .D(SRAM_WE_N_1254), 
         .Z(state_7__N_1453[2])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i2_4_lut.init = 16'hecff;
    LUT4 i1_4_lut_adj_669 (.A(SRAM_WE_N_1254), .B(n20_adj_2522), .C(state[3]), 
         .D(n22), .Z(state_7__N_1453[3])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_4_lut_adj_669.init = 16'hfddd;
    LUT4 i6860_4_lut (.A(state[3]), .B(SRAM_WE_N_1254), .C(n4_adj_2521), 
         .D(n11), .Z(state_7__N_1453[5])) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i6860_4_lut.init = 16'hc8c0;
    LUT4 state_4__bdd_4_lut (.A(state[4]), .B(n18260), .C(SRAM_WE_N_1254), 
         .D(n17319), .Z(LOGIC_CLOCK_enable_46)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C (D))+!B))) */ ;
    defparam state_4__bdd_4_lut.init = 16'h0cec;
    LUT4 i13042_2_lut_4_lut_4_lut (.A(n17336), .B(n17319), .C(SRAM_WE_N_1254), 
         .D(state[4]), .Z(LOGIC_CLOCK_enable_213)) /* synthesis lut_function=(!(A+(B (C)+!B (C (D))))) */ ;
    defparam i13042_2_lut_4_lut_4_lut.init = 16'h0515;
    PFUMX i13266 (.BLUT(n17006), .ALUT(n17005), .C0(state[4]), .Z(n17007));
    LUT4 i3808_3_lut (.A(n7159), .B(n7158), .C(n7130), .Z(\lastAddress[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3808_3_lut.init = 16'hcaca;
    LUT4 i3709_3_lut (.A(n7060), .B(n7059), .C(n7058), .Z(\lastAddress[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3709_3_lut.init = 16'hcaca;
    LUT4 i3805_3_lut (.A(n7156), .B(n7155), .C(n7130), .Z(\lastAddress[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3805_3_lut.init = 16'hcaca;
    LUT4 i3741_3_lut (.A(n7092), .B(n7091), .C(n7090), .Z(\lastAddress[9] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3741_3_lut.init = 16'hcaca;
    LUT4 i3769_3_lut (.A(n7120), .B(n7119), .C(n7118), .Z(\lastAddress[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3769_3_lut.init = 16'hcaca;
    LUT4 i7107_3_lut_3_lut (.A(n17345), .B(n17282), .C(n18260), .Z(LOGIC_CLOCK_enable_47)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+!(C)))) */ ;
    defparam i7107_3_lut_3_lut.init = 16'h4747;
    LUT4 i3761_3_lut (.A(n7112), .B(n7111), .C(n7110), .Z(\lastAddress[14] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3761_3_lut.init = 16'hcaca;
    LUT4 i13089_2_lut_4_lut_4_lut (.A(n17345), .B(n17319), .C(SRAM_WE_N_1254), 
         .D(state[4]), .Z(SRAM_WE_N_1245)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i13089_2_lut_4_lut_4_lut.init = 16'h5040;
    LUT4 i3757_3_lut (.A(n7108), .B(n7107), .C(n7106), .Z(\lastAddress[13] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3757_3_lut.init = 16'hcaca;
    LUT4 i3753_3_lut (.A(n7104), .B(n7103), .C(n7102), .Z(\lastAddress[12] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3753_3_lut.init = 16'hcaca;
    CCU2D lastAddress_31__I_0_304_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(lastAddress_31__N_1310), .B1(\lastAddress[31] ), 
          .C1(\BUS_ADDR_INTERNAL[18]_derived_1 ), .D1(lastAddress[18]), 
          .COUT(n13656));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[12:37])
    defparam lastAddress_31__I_0_304_0.INIT0 = 16'hF000;
    defparam lastAddress_31__I_0_304_0.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_304_0.INJECT1_0 = "NO";
    defparam lastAddress_31__I_0_304_0.INJECT1_1 = "YES";
    LUT4 i6910_3_lut_rep_274_4_lut (.A(state[5]), .B(n17356), .C(SRAM_WE_N_1254), 
         .D(state[4]), .Z(n17282)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i6910_3_lut_rep_274_4_lut.init = 16'hf0e0;
    LUT4 state_7__I_180_i5_4_lut_4_lut (.A(n18260), .B(n51_adj_2510), .C(SRAM_WE_N_1254), 
         .D(n17346), .Z(state_7__N_1453[4])) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B+!(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam state_7__I_180_i5_4_lut_4_lut.init = 16'hc5f5;
    LUT4 i5_4_lut_4_lut (.A(n18260), .B(n17287), .C(n7), .D(n9), .Z(n6250)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i5_4_lut_4_lut.init = 16'h4000;
    LUT4 i6912_2_lut_4_lut_3_lut_4_lut (.A(state[5]), .B(n17356), .C(SRAM_WE_N_1254), 
         .D(state[4]), .Z(SRAM_OE_N_1511)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i6912_2_lut_4_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_311_3_lut_4_lut (.A(state[0]), .B(n17440), .C(state[5]), 
         .D(state[3]), .Z(n17319)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i1_2_lut_rep_311_3_lut_4_lut.init = 16'hfffe;
    CCU2D lastAddress_31__I_0_304_25 (.A0(n17325), .B0(\lastAddress[9] ), 
          .C0(n17337), .D0(\lastAddress[8] ), .A1(n17334), .B1(\lastAddress[7] ), 
          .C1(n17321), .D1(lastAddress[6]), .CIN(n13658), .COUT(n13659));
    defparam lastAddress_31__I_0_304_25.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_304_25.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_304_25.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_304_25.INJECT1_1 = "YES";
    LUT4 i3765_3_lut (.A(n7116), .B(n7115), .C(n7114), .Z(\lastAddress[15] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3765_3_lut.init = 16'hcaca;
    LUT4 lastAddress_i1_i12_3_lut (.A(lastAddress_c[11]), .B(\BUS_addr[11] ), 
         .C(SRAM_WE_N_1254), .Z(n66_c[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam lastAddress_i1_i12_3_lut.init = 16'hacac;
    LUT4 i3749_3_lut (.A(n7100), .B(n7099), .C(n7098), .Z(lastAddress_c[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3749_3_lut.init = 16'hcaca;
    LUT4 i53_4_lut (.A(state[3]), .B(n5990), .C(state[0]), .D(n17440), 
         .Z(n49_adj_2509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i53_4_lut.init = 16'hcfca;
    LUT4 i1_3_lut_4_lut_adj_670 (.A(state[1]), .B(n17455), .C(state[2]), 
         .D(state[3]), .Z(n20)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_670.init = 16'h00f1;
    LUT4 i1_3_lut_4_lut_adj_671 (.A(state[1]), .B(n17455), .C(state[3]), 
         .D(state[2]), .Z(n20_adj_2522)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_671.init = 16'h00f1;
    LUT4 i3737_3_lut (.A(n7088), .B(n7087), .C(n7086), .Z(\lastAddress[8] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i3737_3_lut.init = 16'hcaca;
    LUT4 state_7__I_180_i1_3_lut (.A(n18260), .B(state_7__N_1461[0]), .C(SRAM_WE_N_1254), 
         .Z(state_7__N_1453[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam state_7__I_180_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_672 (.A(state[5]), .B(state[0]), .C(n17007), .D(n5990), 
         .Z(state_7__N_1461[0])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[4] 109[11])
    defparam i1_4_lut_adj_672.init = 16'hdc50;
    
endmodule
//
// Verilog Description of module MatrixDriver
//

module MatrixDriver (MATRIX_CURRROW, PIXEL_CLOCK, PIXEL_CLOCK_N_293, WRITE_DONE, 
            LOGIC_CLOCK_N_57, n18280, currPWMCount, LOGIC_CLOCK, Matrix_CTRL_Out_c_1, 
            currPixel, GND_net, Matrix_LINE_SEL_Out_c_1, n17305, n17380, 
            n13509, n15436, n17278, n17373, n18260, \currPWMCountMax[1] , 
            \currPWMCountMax[2] , \currPWMCountMax[3] , \currPWMCountMax[4] , 
            \currPWMCountMax[5] , \currPWMCountMax[6] , LOGIC_CLOCK_N_57_enable_6, 
            \BUS_data[3] , \currPWMCountMax[10] , \currPWMCountMax[12] , 
            \PWMArray[0][9] , \currPWMCountMax[0] , Matrix_LINE_SEL_Out_c_0, 
            n17411, n17458, n16456, n17368, \SpriteRead_yValid_N_1158[4] , 
            n8, n17371, n17382, n17374, n17329, \currPWMCount[12] , 
            \currPWMCount[11] , \currPWMCount[6] , \currPWMCount[5] , 
            \currPWMCount[4] , \currPWMCount[3] , \currPWMCount[2] , \currPWMCount[1] , 
            \BUS_data[2] , \BUS_data[0] , \BUS_data[1] , \currPWMCountMax[11] , 
            \currPWMCountMax[9] , \currPWMCountMax[8] , \currPWMCountMax[7] , 
            n17326, n17366, n17407, n17453, n17452, \SpriteRead_yValid_N_1158[2] , 
            n15549, n17289, n17408, \SpriteRead_yValid_N_1158[1] , \SpriteRead_yValid_N_1158[0] , 
            n4, Matrix_CTRL_Out_c_2, n15705, n1840, \BUS_currGrantID[0] , 
            \BUS_currGrantID[1] , \BUS_ADDR_INTERNAL[18] , lastAddress_31__N_1310, 
            \BUS_ADDR_INTERNAL[16] , n18277, \BUS_ADDR_INTERNAL[17] , 
            n18264, \BUS_ADDR_INTERNAL[14] , n18262, \BUS_ADDR_INTERNAL[15] , 
            n18271, n3296, Matrix_DATA_Out_c_11, Matrix_DATA_Out_c_10, 
            Matrix_DATA_Out_c_9, Matrix_DATA_Out_c_8, Matrix_DATA_Out_c_7, 
            Matrix_DATA_Out_c_6, Matrix_DATA_Out_c_5, \BUS_ADDR_INTERNAL[12] , 
            n18272, \BUS_ADDR_INTERNAL[13] , n18266, Matrix_DATA_Out_c_4, 
            Matrix_DATA_Out_c_3, Matrix_DATA_Out_c_2, \BUS_ADDR_INTERNAL[10] , 
            n18269, \BUS_ADDR_INTERNAL[11] , n18273, \BUS_ADDR_INTERNAL[8] , 
            n18267, \BUS_ADDR_INTERNAL[9] , n18268, \BUS_ADDR_INTERNAL[7] , 
            n18274, Matrix_DATA_Out_c_1, Matrix_DATA_Out_c_0, Matrix_LINE_SEL_Out_c_2, 
            Matrix_CTRL_Out_c_0, \SpriteRead_yValid_N_1158[3] , n17299, 
            \BUS_ADDR_INTERNAL[5] , n18265, \BUS_ADDR_INTERNAL[6] , n18276, 
            \BUS_ADDR_INTERNAL[3] , n17409, \BUS_ADDR_INTERNAL[4] , n18275, 
            \BUS_ADDR_INTERNAL[1] , n17423, \BUS_ADDR_INTERNAL[2] , n18263, 
            \BUS_ADDR_INTERNAL[0] , n18261, \SpriteRead_yInSprite_7__N_597[0] , 
            n17328, n15539, n17304, n161, n160, n159, n15633, 
            n17307, VRAM_DATA, \VRAM_ADDR[8] , \VRAM_ADDR[7] , \VRAM_ADDR[6] , 
            \VRAM_ADDR[5] , \VRAM_ADDR[4] , \VRAM_ADDR[3] , \VRAM_ADDR[2] , 
            \VRAM_ADDR[1] , \VRAM_ADDR[0] , VRAM_WC, VCC_net, VRAM_WE, 
            VRAM_DATA_OUT);
    output [4:0]MATRIX_CURRROW;
    input PIXEL_CLOCK;
    input PIXEL_CLOCK_N_293;
    output WRITE_DONE;
    input LOGIC_CLOCK_N_57;
    input n18280;
    output [15:0]currPWMCount;
    input LOGIC_CLOCK;
    output Matrix_CTRL_Out_c_1;
    output [7:0]currPixel;
    input GND_net;
    output Matrix_LINE_SEL_Out_c_1;
    input n17305;
    input n17380;
    output n13509;
    input n15436;
    output n17278;
    input n17373;
    input n18260;
    output \currPWMCountMax[1] ;
    output \currPWMCountMax[2] ;
    output \currPWMCountMax[3] ;
    output \currPWMCountMax[4] ;
    output \currPWMCountMax[5] ;
    output \currPWMCountMax[6] ;
    input LOGIC_CLOCK_N_57_enable_6;
    input \BUS_data[3] ;
    output \currPWMCountMax[10] ;
    output \currPWMCountMax[12] ;
    output \PWMArray[0][9] ;
    output \currPWMCountMax[0] ;
    output Matrix_LINE_SEL_Out_c_0;
    input n17411;
    input n17458;
    output n16456;
    output n17368;
    input \SpriteRead_yValid_N_1158[4] ;
    output n8;
    input n17371;
    input n17382;
    input n17374;
    input n17329;
    output \currPWMCount[12] ;
    output \currPWMCount[11] ;
    output \currPWMCount[6] ;
    output \currPWMCount[5] ;
    output \currPWMCount[4] ;
    output \currPWMCount[3] ;
    output \currPWMCount[2] ;
    output \currPWMCount[1] ;
    input \BUS_data[2] ;
    input \BUS_data[0] ;
    input \BUS_data[1] ;
    output \currPWMCountMax[11] ;
    output \currPWMCountMax[9] ;
    output \currPWMCountMax[8] ;
    output \currPWMCountMax[7] ;
    output n17326;
    output n17366;
    output n17407;
    output n17453;
    output n17452;
    input \SpriteRead_yValid_N_1158[2] ;
    output n15549;
    output n17289;
    output n17408;
    input \SpriteRead_yValid_N_1158[1] ;
    input \SpriteRead_yValid_N_1158[0] ;
    output n4;
    output Matrix_CTRL_Out_c_2;
    input n15705;
    input n1840;
    input \BUS_currGrantID[0] ;
    input \BUS_currGrantID[1] ;
    input \BUS_ADDR_INTERNAL[18] ;
    input lastAddress_31__N_1310;
    input \BUS_ADDR_INTERNAL[16] ;
    input n18277;
    input \BUS_ADDR_INTERNAL[17] ;
    input n18264;
    input \BUS_ADDR_INTERNAL[14] ;
    input n18262;
    input \BUS_ADDR_INTERNAL[15] ;
    input n18271;
    input n3296;
    output Matrix_DATA_Out_c_11;
    output Matrix_DATA_Out_c_10;
    output Matrix_DATA_Out_c_9;
    output Matrix_DATA_Out_c_8;
    output Matrix_DATA_Out_c_7;
    output Matrix_DATA_Out_c_6;
    output Matrix_DATA_Out_c_5;
    input \BUS_ADDR_INTERNAL[12] ;
    input n18272;
    input \BUS_ADDR_INTERNAL[13] ;
    input n18266;
    output Matrix_DATA_Out_c_4;
    output Matrix_DATA_Out_c_3;
    output Matrix_DATA_Out_c_2;
    input \BUS_ADDR_INTERNAL[10] ;
    input n18269;
    input \BUS_ADDR_INTERNAL[11] ;
    input n18273;
    input \BUS_ADDR_INTERNAL[8] ;
    input n18267;
    input \BUS_ADDR_INTERNAL[9] ;
    input n18268;
    input \BUS_ADDR_INTERNAL[7] ;
    input n18274;
    output Matrix_DATA_Out_c_1;
    output Matrix_DATA_Out_c_0;
    output Matrix_LINE_SEL_Out_c_2;
    output Matrix_CTRL_Out_c_0;
    input \SpriteRead_yValid_N_1158[3] ;
    output n17299;
    input \BUS_ADDR_INTERNAL[5] ;
    input n18265;
    input \BUS_ADDR_INTERNAL[6] ;
    input n18276;
    input \BUS_ADDR_INTERNAL[3] ;
    input n17409;
    input \BUS_ADDR_INTERNAL[4] ;
    input n18275;
    input \BUS_ADDR_INTERNAL[1] ;
    input n17423;
    input \BUS_ADDR_INTERNAL[2] ;
    input n18263;
    input \BUS_ADDR_INTERNAL[0] ;
    input n18261;
    output \SpriteRead_yInSprite_7__N_597[0] ;
    input n17328;
    input n15539;
    output n17304;
    output n161;
    output n160;
    output n159;
    input n15633;
    output n17307;
    input [29:0]VRAM_DATA;
    input \VRAM_ADDR[8] ;
    input \VRAM_ADDR[7] ;
    input \VRAM_ADDR[6] ;
    input \VRAM_ADDR[5] ;
    input \VRAM_ADDR[4] ;
    input \VRAM_ADDR[3] ;
    input \VRAM_ADDR[2] ;
    input \VRAM_ADDR[1] ;
    input \VRAM_ADDR[0] ;
    input VRAM_WC;
    input VCC_net;
    input VRAM_WE;
    output [29:0]VRAM_DATA_OUT;
    
    wire PIXEL_CLOCK /* synthesis SET_AS_NETWORK=PIXEL_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(43[8:19])
    wire PIXEL_CLOCK_N_293 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(88[9:22])
    wire LOGIC_CLOCK_N_57 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(91[8:15])
    wire [4:0]n12;
    wire [3:0]currBit;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    
    wire PIXEL_CLOCK_enable_9, PIXEL_CLOCK_enable_13;
    wire [3:0]n21;
    
    wire MATRIX_CLKEN_LAT, MATRIX_CLKEN, n15843, n15844, n15847, PWMArray_0__12__N_107, 
        LOGIC_CLOCK_enable_69;
    wire [15:0]currPWMCount_15__N_146;
    
    wire n15845, n15846, n15848, PIXEL_CLOCK_enable_3, n14612, n3, 
        n15850, n15851, n15854, n15852, n15853, n15855, n15773, 
        n15774, n15777, n14157;
    wire [7:0]n37;
    
    wire PIXEL_CLOCK_enable_5, n17354, n14156, n17438, n8_c, n15572, 
        n14155, PIXEL_CLOCK_N_293_enable_26, n7196, n17437, n7187, 
        n7, n14007;
    wire [15:0]currPWMCount_15__N_254;
    
    wire n14008, n17436, n7_adj_2485;
    wire [15:0]currPWMCountMax_15__N_222;
    
    wire n17492, n17493;
    wire [15:0]currPWMVal_15__N_205;
    wire [9:0]\BLUE[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(76[9:13])
    
    wire n15837, n15836, n14006;
    wire [9:0]\RED[1] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(74[9:12])
    
    wire n15832, n15831, n15775, n15776, n15778;
    wire [15:0]\PWMArray[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(79[9:17])
    
    wire n15830, n15829;
    wire [9:0]\GREEN[1] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(75[9:14])
    
    wire n15825;
    wire [15:0]currPWMVal;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(91[9:19])
    
    wire n14154, n15824, n15823, n7191, n5084, n15822;
    wire [9:0]\BLUE[1] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(76[9:13])
    
    wire n15818, n15817, n15816, n15815;
    wire [9:0]\RED[2] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(74[9:12])
    
    wire n15811, n15810, n15809, n15808;
    wire [9:0]\GREEN[2] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(75[9:14])
    
    wire n15804, n15803, n15802, n15801;
    wire [9:0]\BLUE[2] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(76[9:13])
    
    wire n15797, PIXEL_CLOCK_enable_7, n17463, n15796, n7190, n115, 
        n15795, n15794, n70, n13454, n17435, n13461, n4_c;
    wire [9:0]\RED[3] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(74[9:12])
    
    wire n15790, n15789, n15780, n15781, n15784, n13489, n13491, 
        n7_adj_2486;
    wire [9:0]\GREEN[3] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(75[9:14])
    
    wire n15782, n15591, n17391, n148, n7_adj_2487, n17467, BUS_VALID_N_110, 
        n2469, n10348, n15, n17464, n17462, PIXEL_CLOCK_enable_8, 
        MATRIX_ROWCLK_N_279, n138, n6;
    wire [15:0]currPWMCount_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(92[9:21])
    
    wire n3_adj_2489, n3_adj_2490, n17486, n17487, n7_adj_2491, n17351;
    wire [7:0]VRAM_READ_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(85[9:23])
    
    wire VRAM_READ_ADDR_7__N_124, n14005, n17478, n14004, n17477, 
        n15783, n15785, n14009, n14010, PIXEL_CLOCK_enable_20;
    wire [7:0]n47;
    
    wire n25, n14003, n28, n22_adj_2493, n30, n26, n17392, n16803, 
        n14096, n4_adj_2494, n14095, n14094, n14093, n14092, n14257, 
        n14091, n14256, n14090, n14255, n14089, n14254, n15779, 
        n8_adj_2495;
    wire [9:0]\BLUE[3] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(76[9:13])
    
    wire n15786, n8_adj_2496, n15793, n8_adj_2497, n15800, n8_adj_2498, 
        n15807, n8_adj_2499, n15814, n8_adj_2500, n17365, n15821, 
        n8_adj_2501, n14253, n15828, n8_adj_2502, n15835, n8_adj_2503, 
        n15842, n8_adj_2504, n14252, n14251, n15849, n8_adj_2505;
    wire [9:0]\GREEN[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(75[9:14])
    
    wire n15856, n8_adj_2506;
    wire [9:0]\RED[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(74[9:12])
    
    wire n6_adj_2507, n25_adj_2508, n15474, n17353, n15791, n15792, 
        n15798, n15799, n15805, n15806, n15812, n15813, n15819, 
        n15820, n15826, n15827, n15833, n15834, n15840, n15841, 
        n139, n15367, n17470, n14209, n14208, n14207, n14206, 
        n15359, n14205, n14204, n14203, n14202, n14201, n14200, 
        n14199, n15839, n9, n15788, n15787, n15838;
    
    FD1S3AX currRow_i0_i0 (.D(n12[0]), .CK(PIXEL_CLOCK), .Q(MATRIX_CURRROW[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam currRow_i0_i0.GSR = "DISABLED";
    FD1P3IX currBit_997__i3 (.D(n21[3]), .SP(PIXEL_CLOCK_enable_9), .CD(PIXEL_CLOCK_enable_13), 
            .CK(PIXEL_CLOCK), .Q(currBit[3]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_997__i3.GSR = "DISABLED";
    FD1S3AX MATRIX_CLKEN_LAT_155 (.D(MATRIX_CLKEN), .CK(PIXEL_CLOCK_N_293), 
            .Q(MATRIX_CLKEN_LAT)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam MATRIX_CLKEN_LAT_155.GSR = "DISABLED";
    PFUMX i12185 (.BLUT(n15843), .ALUT(n15844), .C0(currBit[1]), .Z(n15847));
    FD1P3IX currBit_997__i2 (.D(n21[2]), .SP(PIXEL_CLOCK_enable_9), .CD(PIXEL_CLOCK_enable_13), 
            .CK(PIXEL_CLOCK), .Q(currBit[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_997__i2.GSR = "DISABLED";
    FD1S3DX WRITE_DONE_158 (.D(n18280), .CK(LOGIC_CLOCK_N_57), .CD(PWMArray_0__12__N_107), 
            .Q(WRITE_DONE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam WRITE_DONE_158.GSR = "DISABLED";
    FD1P3BX currPWMCount_i0 (.D(currPWMCount_15__N_146[0]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i0.GSR = "DISABLED";
    PFUMX i12186 (.BLUT(n15845), .ALUT(n15846), .C0(currBit[1]), .Z(n15848));
    FD1P3IX MATRIX_CLKEN_145 (.D(n18280), .SP(PIXEL_CLOCK_enable_3), .CD(n14612), 
            .CK(PIXEL_CLOCK), .Q(MATRIX_CLKEN)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam MATRIX_CLKEN_145.GSR = "DISABLED";
    FD1P3IX currBit_997__i1 (.D(n3), .SP(PIXEL_CLOCK_enable_9), .CD(PIXEL_CLOCK_enable_13), 
            .CK(PIXEL_CLOCK), .Q(currBit[1]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_997__i1.GSR = "DISABLED";
    PFUMX i12192 (.BLUT(n15850), .ALUT(n15851), .C0(currBit[1]), .Z(n15854));
    PFUMX i12193 (.BLUT(n15852), .ALUT(n15853), .C0(currBit[1]), .Z(n15855));
    PFUMX i12115 (.BLUT(n15773), .ALUT(n15774), .C0(currBit[1]), .Z(n15777));
    CCU2D currPixel_996_add_4_9 (.A0(currPixel[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14157), .S0(n37[7]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_add_4_9.INIT0 = 16'hfaaa;
    defparam currPixel_996_add_4_9.INIT1 = 16'h0000;
    defparam currPixel_996_add_4_9.INJECT1_0 = "NO";
    defparam currPixel_996_add_4_9.INJECT1_1 = "NO";
    FD1P3AX MATRIX_ROWLAT_149 (.D(n17354), .SP(PIXEL_CLOCK_enable_5), .CK(PIXEL_CLOCK), 
            .Q(Matrix_LINE_SEL_Out_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam MATRIX_ROWLAT_149.GSR = "DISABLED";
    CCU2D currPixel_996_add_4_7 (.A0(currPixel[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14156), .COUT(n14157), .S0(n37[5]), .S1(n37[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_add_4_7.INIT0 = 16'hfaaa;
    defparam currPixel_996_add_4_7.INIT1 = 16'hfaaa;
    defparam currPixel_996_add_4_7.INJECT1_0 = "NO";
    defparam currPixel_996_add_4_7.INJECT1_1 = "NO";
    FD1P3IX currBit_997__i0 (.D(n17438), .SP(PIXEL_CLOCK_enable_9), .CD(PIXEL_CLOCK_enable_13), 
            .CK(PIXEL_CLOCK), .Q(currBit[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_997__i0.GSR = "DISABLED";
    LUT4 i4_4_lut (.A(n17305), .B(n8_c), .C(n17380), .D(n15572), .Z(n13509)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i3_4_lut (.A(n15436), .B(n17278), .C(n17373), .D(n18260), .Z(n8_c)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    CCU2D currPixel_996_add_4_5 (.A0(currPixel[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14155), .COUT(n14156), .S0(n37[3]), .S1(n37[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_add_4_5.INIT0 = 16'hfaaa;
    defparam currPixel_996_add_4_5.INIT1 = 16'hfaaa;
    defparam currPixel_996_add_4_5.INJECT1_0 = "NO";
    defparam currPixel_996_add_4_5.INJECT1_1 = "NO";
    FD1P3IX currPWMCountMax__i2 (.D(n3), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7196), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i2.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i3 (.D(n17437), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7196), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i3.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i4 (.D(n7), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i4.GSR = "DISABLED";
    CCU2D add_107_11 (.A0(currPWMCount[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14007), .COUT(n14008), .S0(currPWMCount_15__N_254[9]), 
          .S1(currPWMCount_15__N_254[10]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_11.INIT0 = 16'h5aaa;
    defparam add_107_11.INIT1 = 16'h5aaa;
    defparam add_107_11.INJECT1_0 = "NO";
    defparam add_107_11.INJECT1_1 = "NO";
    FD1P3IX currPWMCountMax__i5 (.D(n17436), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i5.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i6 (.D(n7_adj_2485), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i6.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .D(currBit[0]), .Z(currPWMCountMax_15__N_222[7])) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B ((D)+!C)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0c18;
    PFUMX i13422 (.BLUT(n17492), .ALUT(n17493), .C0(currBit[0]), .Z(currPWMVal_15__N_205[11]));
    LUT4 i12175_3_lut (.A(\BLUE[0] [2]), .B(\BLUE[0] [3]), .C(currBit[0]), 
         .Z(n15837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12175_3_lut.init = 16'hcaca;
    LUT4 i12174_3_lut (.A(\BLUE[0] [0]), .B(\BLUE[0] [1]), .C(currBit[0]), 
         .Z(n15836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12174_3_lut.init = 16'hcaca;
    CCU2D add_107_9 (.A0(currPWMCount[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14006), .COUT(n14007), .S0(currPWMCount_15__N_254[7]), 
          .S1(currPWMCount_15__N_254[8]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_9.INIT0 = 16'h5aaa;
    defparam add_107_9.INIT1 = 16'h5aaa;
    defparam add_107_9.INJECT1_0 = "NO";
    defparam add_107_9.INJECT1_1 = "NO";
    LUT4 i12170_3_lut (.A(\RED[1] [6]), .B(\RED[1] [7]), .C(currBit[0]), 
         .Z(n15832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12170_3_lut.init = 16'hcaca;
    LUT4 i12169_3_lut (.A(\RED[1] [4]), .B(\RED[1] [5]), .C(currBit[0]), 
         .Z(n15831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12169_3_lut.init = 16'hcaca;
    PFUMX i12116 (.BLUT(n15775), .ALUT(n15776), .C0(currBit[1]), .Z(n15778));
    FD1P3IX currPWMCountMax__i7 (.D(currBit[2]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i7.GSR = "DISABLED";
    FD1P3AY brightness_3__159 (.D(\BUS_data[3] ), .SP(LOGIC_CLOCK_N_57_enable_6), 
            .CK(LOGIC_CLOCK_N_57), .Q(\PWMArray[0] [12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam brightness_3__159.GSR = "DISABLED";
    LUT4 i12168_3_lut (.A(\RED[1] [2]), .B(\RED[1] [3]), .C(currBit[0]), 
         .Z(n15830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12168_3_lut.init = 16'hcaca;
    LUT4 i12167_3_lut (.A(\RED[1] [0]), .B(\RED[1] [1]), .C(currBit[0]), 
         .Z(n15829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12167_3_lut.init = 16'hcaca;
    LUT4 i12163_3_lut (.A(\GREEN[1] [6]), .B(\GREEN[1] [7]), .C(currBit[0]), 
         .Z(n15825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12163_3_lut.init = 16'hcaca;
    FD1P3AX currPWMVal_i0_i11 (.D(currPWMVal_15__N_205[11]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i11.GSR = "DISABLED";
    CCU2D currPixel_996_add_4_3 (.A0(currPixel[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14154), .COUT(n14155), .S0(n37[1]), .S1(n37[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_add_4_3.INIT0 = 16'hfaaa;
    defparam currPixel_996_add_4_3.INIT1 = 16'hfaaa;
    defparam currPixel_996_add_4_3.INJECT1_0 = "NO";
    defparam currPixel_996_add_4_3.INJECT1_1 = "NO";
    LUT4 i12162_3_lut (.A(\GREEN[1] [4]), .B(\GREEN[1] [5]), .C(currBit[0]), 
         .Z(n15824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12162_3_lut.init = 16'hcaca;
    LUT4 i12161_3_lut (.A(\GREEN[1] [2]), .B(\GREEN[1] [3]), .C(currBit[0]), 
         .Z(n15823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12161_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[0]), 
         .D(currBit[3]), .Z(currPWMCountMax_15__N_222[9])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B+!((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i22_4_lut_4_lut.init = 16'h1181;
    FD1P3AX currPWMVal_i0_i10 (.D(currPWMVal_15__N_205[10]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i10.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i11 (.D(n5084), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7191), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i11.GSR = "DISABLED";
    LUT4 i12160_3_lut (.A(\GREEN[1] [0]), .B(\GREEN[1] [1]), .C(currBit[0]), 
         .Z(n15822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12160_3_lut.init = 16'hcaca;
    LUT4 i12156_3_lut (.A(\BLUE[1] [6]), .B(\BLUE[1] [7]), .C(currBit[0]), 
         .Z(n15818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12156_3_lut.init = 16'hcaca;
    LUT4 i12155_3_lut (.A(\BLUE[1] [4]), .B(\BLUE[1] [5]), .C(currBit[0]), 
         .Z(n15817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12155_3_lut.init = 16'hcaca;
    FD1P3AX currPWMVal_i0_i9 (.D(currPWMVal_15__N_205[9]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i9.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i8 (.D(currPWMVal_15__N_205[8]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i8.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i7 (.D(currPWMVal_15__N_205[7]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i7.GSR = "DISABLED";
    LUT4 i12154_3_lut (.A(\BLUE[1] [2]), .B(\BLUE[1] [3]), .C(currBit[0]), 
         .Z(n15816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12154_3_lut.init = 16'hcaca;
    LUT4 i12153_3_lut (.A(\BLUE[1] [0]), .B(\BLUE[1] [1]), .C(currBit[0]), 
         .Z(n15815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12153_3_lut.init = 16'hcaca;
    CCU2D currPixel_996_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n14154), .S1(n37[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_add_4_1.INIT0 = 16'hF000;
    defparam currPixel_996_add_4_1.INIT1 = 16'h0555;
    defparam currPixel_996_add_4_1.INJECT1_0 = "NO";
    defparam currPixel_996_add_4_1.INJECT1_1 = "NO";
    LUT4 i12149_3_lut (.A(\RED[2] [6]), .B(\RED[2] [7]), .C(currBit[0]), 
         .Z(n15811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12149_3_lut.init = 16'hcaca;
    LUT4 i12148_3_lut (.A(\RED[2] [4]), .B(\RED[2] [5]), .C(currBit[0]), 
         .Z(n15810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12148_3_lut.init = 16'hcaca;
    LUT4 i12147_3_lut (.A(\RED[2] [2]), .B(\RED[2] [3]), .C(currBit[0]), 
         .Z(n15809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12147_3_lut.init = 16'hcaca;
    LUT4 i12146_3_lut (.A(\RED[2] [0]), .B(\RED[2] [1]), .C(currBit[0]), 
         .Z(n15808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12146_3_lut.init = 16'hcaca;
    LUT4 i12142_3_lut (.A(\GREEN[2] [6]), .B(\GREEN[2] [7]), .C(currBit[0]), 
         .Z(n15804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12142_3_lut.init = 16'hcaca;
    LUT4 i12141_3_lut (.A(\GREEN[2] [4]), .B(\GREEN[2] [5]), .C(currBit[0]), 
         .Z(n15803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12141_3_lut.init = 16'hcaca;
    LUT4 i12140_3_lut (.A(\GREEN[2] [2]), .B(\GREEN[2] [3]), .C(currBit[0]), 
         .Z(n15802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12140_3_lut.init = 16'hcaca;
    LUT4 i12139_3_lut (.A(\GREEN[2] [0]), .B(\GREEN[2] [1]), .C(currBit[0]), 
         .Z(n15801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12139_3_lut.init = 16'hcaca;
    LUT4 i12135_3_lut (.A(\BLUE[2] [6]), .B(\BLUE[2] [7]), .C(currBit[0]), 
         .Z(n15797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12135_3_lut.init = 16'hcaca;
    FD1P3AX MATRIX_LAT_146 (.D(n17463), .SP(PIXEL_CLOCK_enable_7), .CK(PIXEL_CLOCK), 
            .Q(Matrix_CTRL_Out_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam MATRIX_LAT_146.GSR = "DISABLED";
    LUT4 i12134_3_lut (.A(\BLUE[2] [4]), .B(\BLUE[2] [5]), .C(currBit[0]), 
         .Z(n15796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12134_3_lut.init = 16'hcaca;
    FD1P3IX currPWMCountMax__i13 (.D(n115), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7190), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i13.GSR = "DISABLED";
    LUT4 i12133_3_lut (.A(\BLUE[2] [2]), .B(\BLUE[2] [3]), .C(currBit[0]), 
         .Z(n15795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12133_3_lut.init = 16'hcaca;
    LUT4 i12132_3_lut (.A(\BLUE[2] [0]), .B(\BLUE[2] [1]), .C(currBit[0]), 
         .Z(n15794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12132_3_lut.init = 16'hcaca;
    LUT4 i10327_4_lut (.A(n70), .B(n13454), .C(currBit[0]), .D(n17435), 
         .Z(currPWMVal_15__N_205[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10327_4_lut.init = 16'hcac0;
    LUT4 i10326_3_lut (.A(\PWMArray[0][9] ), .B(\PWMArray[0] [11]), .C(currBit[3]), 
         .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10326_3_lut.init = 16'hcaca;
    LUT4 i10310_3_lut (.A(n13454), .B(n13461), .C(currBit[0]), .Z(currPWMVal_15__N_205[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10310_3_lut.init = 16'hcaca;
    LUT4 i10332_4_lut (.A(n13461), .B(currBit[2]), .C(currBit[0]), .D(n4_c), 
         .Z(currPWMVal_15__N_205[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10332_4_lut.init = 16'hca0a;
    LUT4 i12128_3_lut (.A(\RED[3] [6]), .B(\RED[3] [7]), .C(currBit[0]), 
         .Z(n15790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12128_3_lut.init = 16'hcaca;
    LUT4 i12127_3_lut (.A(\RED[3] [4]), .B(\RED[3] [5]), .C(currBit[0]), 
         .Z(n15789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12127_3_lut.init = 16'hcaca;
    PFUMX i12122 (.BLUT(n15780), .ALUT(n15781), .C0(currBit[1]), .Z(n15784));
    LUT4 i2_3_lut_4_lut (.A(\PWMArray[0][9] ), .B(n17435), .C(currBit[0]), 
         .D(currBit[3]), .Z(currPWMVal_15__N_205[0])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 i10350_3_lut (.A(n13489), .B(n13491), .C(currBit[0]), .Z(n7_adj_2486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10350_3_lut.init = 16'hcaca;
    LUT4 i10572_3_lut_4_lut (.A(currBit[1]), .B(currBit[0]), .C(currBit[2]), 
         .D(currBit[3]), .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10572_3_lut_4_lut.init = 16'h7f80;
    LUT4 i10565_2_lut_3_lut (.A(currBit[1]), .B(currBit[0]), .C(currBit[2]), 
         .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10565_2_lut_3_lut.init = 16'h7878;
    FD1P3IX currPWMVal_i0_i4 (.D(n7_adj_2486), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i4.GSR = "DISABLED";
    LUT4 i12120_3_lut (.A(\GREEN[3] [4]), .B(\GREEN[3] [5]), .C(currBit[0]), 
         .Z(n15782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12120_3_lut.init = 16'hcaca;
    LUT4 i13121_2_lut_rep_427 (.A(currBit[1]), .B(currBit[2]), .Z(n17435)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i13121_2_lut_rep_427.init = 16'h1111;
    LUT4 i11936_2_lut_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .D(currBit[0]), .Z(n15591)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11936_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i13113_2_lut_3_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .Z(n115)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i13113_2_lut_3_lut.init = 16'h0101;
    LUT4 i6771_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .D(currBit[0]), .Z(currPWMCountMax_15__N_222[11])) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;
    defparam i6771_3_lut_4_lut.init = 16'h1001;
    LUT4 i1_2_lut_rep_383_3_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[0]), 
         .Z(n17391)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_383_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(currBit[1]), .B(currBit[2]), .C(\PWMArray[0] [10]), 
         .Z(n148)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    FD1P3IX currPWMVal_i0_i5 (.D(n7_adj_2487), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i5.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i6 (.D(currPWMVal_15__N_205[6]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i6.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i12 (.D(currPWMVal_15__N_205[12]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i12.GSR = "DISABLED";
    LUT4 i809_2_lut_rep_428 (.A(currBit[1]), .B(currBit[2]), .Z(n17436)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(195[36:65])
    defparam i809_2_lut_rep_428.init = 16'h6666;
    LUT4 i10424_3_lut_3_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[0]), 
         .Z(n7)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(195[36:65])
    defparam i10424_3_lut_3_lut.init = 16'h3636;
    LUT4 i10422_3_lut_3_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[0]), 
         .Z(n7_adj_2485)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(195[36:65])
    defparam i10422_3_lut_3_lut.init = 16'h6c6c;
    LUT4 i12006_2_lut_rep_429 (.A(currBit[0]), .B(currBit[1]), .Z(n17437)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12006_2_lut_rep_429.init = 16'heeee;
    LUT4 i3_3_lut_4_lut (.A(currBit[0]), .B(currBit[1]), .C(currBit[3]), 
         .D(n17467), .Z(currPWMVal_15__N_205[12])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0100;
    LUT4 i10556_1_lut_rep_430 (.A(currBit[0]), .Z(n17438)) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10556_1_lut_rep_430.init = 16'h5555;
    LUT4 i1_3_lut_3_lut (.A(currBit[0]), .B(currBit[3]), .C(currBit[1]), 
         .Z(n5084)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_3_lut_3_lut.init = 16'h0d0d;
    LUT4 BUS_VALID_I_7_2_lut_rep_270 (.A(BUS_VALID_N_110), .B(n2469), .Z(n17278)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(269[29:83])
    defparam BUS_VALID_I_7_2_lut_rep_270.init = 16'h2222;
    FD1P3IX currPWMCountMax__i1 (.D(n115), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n10348), .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i1.GSR = "DISABLED";
    LUT4 i10338_4_lut (.A(currBit[2]), .B(n13489), .C(currBit[0]), .D(n15), 
         .Z(n7_adj_2487)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10338_4_lut.init = 16'hcac0;
    LUT4 i10334_3_lut (.A(\PWMArray[0] [11]), .B(\PWMArray[0][9] ), .C(currBit[1]), 
         .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10334_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n17464), .B(n17462), .C(n15), .D(currBit[0]), 
         .Z(currPWMVal_15__N_205[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i1_4_lut.init = 16'hc088;
    FD1P3AX MATRIX_ROWCLK_148 (.D(MATRIX_ROWCLK_N_279), .SP(PIXEL_CLOCK_enable_8), 
            .CK(PIXEL_CLOCK), .Q(Matrix_LINE_SEL_Out_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam MATRIX_ROWCLK_148.GSR = "DISABLED";
    LUT4 PWMArray_0__12__I_6_2_lut_3_lut (.A(BUS_VALID_N_110), .B(n2469), 
         .C(n18260), .Z(PWMArray_0__12__N_107)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(269[29:83])
    defparam PWMArray_0__12__I_6_2_lut_3_lut.init = 16'hfdfd;
    LUT4 i13073_3_lut_4_lut (.A(BUS_VALID_N_110), .B(n2469), .C(n17411), 
         .D(n17458), .Z(n16456)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(269[29:83])
    defparam i13073_3_lut_4_lut.init = 16'hd000;
    LUT4 i1_4_lut_4_lut (.A(currBit[2]), .B(currBit[3]), .C(\PWMArray[0] [12]), 
         .D(\PWMArray[0] [10]), .Z(n138)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_4_lut_4_lut.init = 16'h5140;
    LUT4 SpriteRead_yInSprite_7__N_597_7__I_0_i8_3_lut_3_lut_4_lut (.A(MATRIX_CURRROW[4]), 
         .B(n17368), .C(n6), .D(\SpriteRead_yValid_N_1158[4] ), .Z(n8)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (B (C (D))+!B (C+(D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam SpriteRead_yInSprite_7__N_597_7__I_0_i8_3_lut_3_lut_4_lut.init = 16'hf990;
    LUT4 i11918_2_lut_3_lut_4_lut (.A(n17371), .B(n17382), .C(n17374), 
         .D(n17329), .Z(n15572)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(275[55:66])
    defparam i11918_2_lut_3_lut_4_lut.init = 16'hfffe;
    FD1P3BX currPWMCount_i15 (.D(currPWMCount_15__N_146[15]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount_c[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i15.GSR = "DISABLED";
    FD1P3BX currPWMCount_i14 (.D(currPWMCount_15__N_146[14]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount_c[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i14.GSR = "DISABLED";
    FD1P3BX currPWMCount_i13 (.D(currPWMCount_15__N_146[13]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount_c[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i13.GSR = "DISABLED";
    FD1P3BX currPWMCount_i12 (.D(currPWMCount_15__N_146[12]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i12.GSR = "DISABLED";
    FD1P3BX currPWMCount_i11 (.D(currPWMCount_15__N_146[11]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i11.GSR = "DISABLED";
    FD1P3BX currPWMCount_i10 (.D(currPWMCount_15__N_146[10]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i10.GSR = "DISABLED";
    FD1P3BX currPWMCount_i9 (.D(currPWMCount_15__N_146[9]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i9.GSR = "DISABLED";
    FD1P3BX currPWMCount_i8 (.D(currPWMCount_15__N_146[8]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i8.GSR = "DISABLED";
    FD1P3BX currPWMCount_i7 (.D(currPWMCount_15__N_146[7]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i7.GSR = "DISABLED";
    FD1P3BX currPWMCount_i6 (.D(currPWMCount_15__N_146[6]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i6.GSR = "DISABLED";
    FD1P3BX currPWMCount_i5 (.D(currPWMCount_15__N_146[5]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i5.GSR = "DISABLED";
    FD1P3BX currPWMCount_i4 (.D(currPWMCount_15__N_146[4]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i4.GSR = "DISABLED";
    FD1P3BX currPWMCount_i3 (.D(currPWMCount_15__N_146[3]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i3.GSR = "DISABLED";
    FD1P3BX currPWMCount_i2 (.D(currPWMCount_15__N_146[2]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i2.GSR = "DISABLED";
    FD1P3BX currPWMCount_i1 (.D(currPWMCount_15__N_146[1]), .SP(LOGIC_CLOCK_enable_69), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(\currPWMCount[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(206[3] 214[10])
    defparam currPWMCount_i1.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i1 (.D(n3_adj_2489), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7196), .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i1.GSR = "DISABLED";
    FD1P3AY brightness_2__160 (.D(\BUS_data[2] ), .SP(LOGIC_CLOCK_N_57_enable_6), 
            .CK(LOGIC_CLOCK_N_57), .Q(\PWMArray[0] [11])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam brightness_2__160.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i2 (.D(n3_adj_2490), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7196), .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i2.GSR = "DISABLED";
    PFUMX i13418 (.BLUT(n17486), .ALUT(n17487), .C0(\PWMArray[0] [11]), 
          .Z(n13461));
    FD1P3IX currPWMVal_i0_i3 (.D(n7_adj_2491), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CD(n7187), .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i3.GSR = "DISABLED";
    FD1P3AY brightness_0__162 (.D(\BUS_data[0] ), .SP(LOGIC_CLOCK_N_57_enable_6), 
            .CK(LOGIC_CLOCK_N_57), .Q(\PWMArray[0][9] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam brightness_0__162.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i0 (.D(currPWMVal_15__N_205[0]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(currPWMVal[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMVal_i0_i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_645 (.A(currPixel[0]), .B(n17351), .C(currPixel[1]), 
         .D(n15591), .Z(PIXEL_CLOCK_enable_8)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C)))) */ ;
    defparam i1_4_lut_adj_645.init = 16'h4048;
    FD1P3AY brightness_1__161 (.D(\BUS_data[1] ), .SP(LOGIC_CLOCK_N_57_enable_6), 
            .CK(LOGIC_CLOCK_N_57), .Q(\PWMArray[0] [10])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam brightness_1__161.GSR = "DISABLED";
    FD1P3AX VRAM_PAGEMAPPING_152 (.D(VRAM_READ_ADDR_7__N_124), .SP(PIXEL_CLOCK_enable_9), 
            .CK(PIXEL_CLOCK), .Q(VRAM_READ_ADDR[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam VRAM_PAGEMAPPING_152.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i12 (.D(currPWMCountMax_15__N_222[11]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i12.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i10 (.D(currPWMCountMax_15__N_222[9]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i10.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i9 (.D(currPWMCountMax_15__N_222[8]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i9.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i8 (.D(currPWMCountMax_15__N_222[7]), .SP(PIXEL_CLOCK_N_293_enable_26), 
            .CK(PIXEL_CLOCK_N_293), .Q(\currPWMCountMax[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(192[3] 198[10])
    defparam currPWMCountMax__i8.GSR = "DISABLED";
    FD1P3AX currRow_i0_i4 (.D(n17326), .SP(PIXEL_CLOCK_enable_13), .CK(PIXEL_CLOCK), 
            .Q(MATRIX_CURRROW[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam currRow_i0_i4.GSR = "DISABLED";
    FD1P3AX currRow_i0_i3 (.D(n17366), .SP(PIXEL_CLOCK_enable_13), .CK(PIXEL_CLOCK), 
            .Q(MATRIX_CURRROW[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam currRow_i0_i3.GSR = "DISABLED";
    FD1P3AX currRow_i0_i2 (.D(n17407), .SP(PIXEL_CLOCK_enable_13), .CK(PIXEL_CLOCK), 
            .Q(MATRIX_CURRROW[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam currRow_i0_i2.GSR = "DISABLED";
    FD1P3AX currRow_i0_i1 (.D(n17453), .SP(PIXEL_CLOCK_enable_13), .CK(PIXEL_CLOCK), 
            .Q(MATRIX_CURRROW[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=142, LSE_RLINE=142 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam currRow_i0_i1.GSR = "DISABLED";
    CCU2D add_107_7 (.A0(\currPWMCount[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[6] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14005), .COUT(n14006), .S0(currPWMCount_15__N_254[5]), 
          .S1(currPWMCount_15__N_254[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_7.INIT0 = 16'h5aaa;
    defparam add_107_7.INIT1 = 16'h5aaa;
    defparam add_107_7.INJECT1_0 = "NO";
    defparam add_107_7.INJECT1_1 = "NO";
    LUT4 i10391_then_4_lut (.A(currBit[0]), .B(currBit[3]), .C(currBit[2]), 
         .D(currBit[1]), .Z(n17478)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i10391_then_4_lut.init = 16'h3337;
    LUT4 i1561_2_lut_rep_444 (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .Z(n17452)) /* synthesis lut_function=(A (B)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1561_2_lut_rep_444.init = 16'h8888;
    LUT4 i1566_2_lut_rep_399_3_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[2]), .Z(n17407)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1566_2_lut_rep_399_3_lut.init = 16'h7878;
    CCU2D add_107_5 (.A0(\currPWMCount[3] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[4] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14004), .COUT(n14005), .S0(currPWMCount_15__N_254[3]), 
          .S1(currPWMCount_15__N_254[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_5.INIT0 = 16'h5aaa;
    defparam add_107_5.INIT1 = 16'h5aaa;
    defparam add_107_5.INJECT1_0 = "NO";
    defparam add_107_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(\SpriteRead_yValid_N_1158[2] ), .D(MATRIX_CURRROW[2]), .Z(n15549)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8778;
    LUT4 i10391_else_4_lut (.A(currBit[0]), .B(currBit[3]), .C(currBit[2]), 
         .D(currBit[1]), .Z(n17477)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i10391_else_4_lut.init = 16'hccc8;
    LUT4 i6746_2_lut (.A(currPWMCount_15__N_254[15]), .B(n17289), .Z(currPWMCount_15__N_146[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6746_2_lut.init = 16'h2222;
    LUT4 i1575_2_lut_rep_360_3_lut_4_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[3]), .D(MATRIX_CURRROW[2]), .Z(n17368)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1575_2_lut_rep_360_3_lut_4_lut.init = 16'h8000;
    LUT4 i1573_2_lut_rep_358_3_lut_4_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[3]), .D(MATRIX_CURRROW[2]), .Z(n17366)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1573_2_lut_rep_358_3_lut_4_lut.init = 16'h78f0;
    LUT4 i6747_2_lut (.A(currPWMCount_15__N_254[14]), .B(n17289), .Z(currPWMCount_15__N_146[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6747_2_lut.init = 16'h2222;
    LUT4 i1568_2_lut_rep_400_3_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[2]), .Z(n17408)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1568_2_lut_rep_400_3_lut.init = 16'h8080;
    LUT4 i6748_2_lut (.A(currPWMCount_15__N_254[13]), .B(n17289), .Z(currPWMCount_15__N_146[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6748_2_lut.init = 16'h2222;
    LUT4 i1559_2_lut_rep_445 (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .Z(n17453)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1559_2_lut_rep_445.init = 16'h6666;
    LUT4 i6749_2_lut (.A(currPWMCount_15__N_254[12]), .B(n17289), .Z(currPWMCount_15__N_146[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6749_2_lut.init = 16'h2222;
    LUT4 SpriteRead_yInSprite_7__N_597_7__I_0_i4_4_lut_4_lut (.A(MATRIX_CURRROW[1]), 
         .B(MATRIX_CURRROW[0]), .C(\SpriteRead_yValid_N_1158[1] ), .D(\SpriteRead_yValid_N_1158[0] ), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C (D))+!B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam SpriteRead_yInSprite_7__N_597_7__I_0_i4_4_lut_4_lut.init = 16'hd890;
    LUT4 i6750_2_lut (.A(currPWMCount_15__N_254[11]), .B(n17289), .Z(currPWMCount_15__N_146[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6750_2_lut.init = 16'h2222;
    LUT4 i6751_2_lut (.A(currPWMCount_15__N_254[10]), .B(n17289), .Z(currPWMCount_15__N_146[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6751_2_lut.init = 16'h2222;
    LUT4 i6752_2_lut (.A(currPWMCount_15__N_254[9]), .B(n17289), .Z(currPWMCount_15__N_146[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6752_2_lut.init = 16'h2222;
    LUT4 i6753_2_lut (.A(currPWMCount_15__N_254[8]), .B(n17289), .Z(currPWMCount_15__N_146[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6753_2_lut.init = 16'h2222;
    LUT4 i6754_2_lut (.A(currPWMCount_15__N_254[7]), .B(n17289), .Z(currPWMCount_15__N_146[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6754_2_lut.init = 16'h2222;
    PFUMX i12123 (.BLUT(n15782), .ALUT(n15783), .C0(currBit[1]), .Z(n15785));
    CCU2D add_107_15 (.A0(currPWMCount_c[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount_c[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14009), .COUT(n14010), .S0(currPWMCount_15__N_254[13]), 
          .S1(currPWMCount_15__N_254[14]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_15.INIT0 = 16'h5aaa;
    defparam add_107_15.INIT1 = 16'h5aaa;
    defparam add_107_15.INJECT1_0 = "NO";
    defparam add_107_15.INJECT1_1 = "NO";
    FD1P3AX currPixel_996__i0 (.D(n47[0]), .SP(PIXEL_CLOCK_enable_20), .CK(PIXEL_CLOCK), 
            .Q(currPixel[0])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i0.GSR = "DISABLED";
    LUT4 i6755_2_lut (.A(currPWMCount_15__N_254[6]), .B(n17289), .Z(currPWMCount_15__N_146[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6755_2_lut.init = 16'h2222;
    CCU2D add_107_17 (.A0(currPWMCount_c[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14010), .S0(currPWMCount_15__N_254[15]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_17.INIT0 = 16'h5aaa;
    defparam add_107_17.INIT1 = 16'h0000;
    defparam add_107_17.INJECT1_0 = "NO";
    defparam add_107_17.INJECT1_1 = "NO";
    LUT4 i6756_2_lut (.A(currPWMCount_15__N_254[5]), .B(n17289), .Z(currPWMCount_15__N_146[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6756_2_lut.init = 16'h2222;
    LUT4 i6757_2_lut (.A(currPWMCount_15__N_254[4]), .B(n17289), .Z(currPWMCount_15__N_146[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6757_2_lut.init = 16'h2222;
    LUT4 i6760_2_lut (.A(currPWMCount_15__N_254[3]), .B(n17289), .Z(currPWMCount_15__N_146[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6760_2_lut.init = 16'h2222;
    LUT4 i6761_2_lut (.A(currPWMCount_15__N_254[2]), .B(n17289), .Z(currPWMCount_15__N_146[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6761_2_lut.init = 16'h2222;
    LUT4 i6762_2_lut (.A(currPWMCount_15__N_254[1]), .B(n17289), .Z(currPWMCount_15__N_146[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6762_2_lut.init = 16'h2222;
    LUT4 i9_4_lut (.A(currPWMCount[0]), .B(\currPWMCount[1] ), .C(\currPWMCount[6] ), 
         .D(\currPWMCount[4] ), .Z(n25)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    CCU2D add_107_3 (.A0(\currPWMCount[1] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[2] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14003), .COUT(n14004), .S0(currPWMCount_15__N_254[1]), 
          .S1(currPWMCount_15__N_254[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_3.INIT0 = 16'h5aaa;
    defparam add_107_3.INIT1 = 16'h5aaa;
    defparam add_107_3.INJECT1_0 = "NO";
    defparam add_107_3.INJECT1_1 = "NO";
    LUT4 i14_4_lut (.A(currPWMCount[10]), .B(n28), .C(n22_adj_2493), .D(\currPWMCount[12] ), 
         .Z(n30)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i14_4_lut.init = 16'h8000;
    LUT4 i10_4_lut (.A(currPWMCount[8]), .B(\currPWMCount[3] ), .C(currPWMCount_c[13]), 
         .D(\currPWMCount[5] ), .Z(n26)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i10_4_lut.init = 16'h8000;
    LUT4 i10415_4_lut (.A(currBit[1]), .B(currBit[0]), .C(\PWMArray[0][9] ), 
         .D(\PWMArray[0] [10]), .Z(n3_adj_2489)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10415_4_lut.init = 16'h6420;
    LUT4 i12_4_lut (.A(\currPWMCount[11] ), .B(currPWMCount[9]), .C(currPWMCount_c[14]), 
         .D(currPWMCount_c[15]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut.init = 16'h8000;
    LUT4 i10383_4_lut (.A(currBit[1]), .B(n15), .C(currBit[0]), .D(\PWMArray[0] [10]), 
         .Z(n3_adj_2490)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10383_4_lut.init = 16'hcac0;
    LUT4 i6_2_lut (.A(\currPWMCount[2] ), .B(currPWMCount[7]), .Z(n22_adj_2493)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6_2_lut.init = 16'h8888;
    LUT4 i10341_4_lut (.A(n13491), .B(currBit[2]), .C(currBit[0]), .D(n17464), 
         .Z(n7_adj_2491)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10341_4_lut.init = 16'h3a0a;
    LUT4 i6567_2_lut (.A(currPWMCount_15__N_254[0]), .B(n17289), .Z(currPWMCount_15__N_146[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(209[4] 213[11])
    defparam i6567_2_lut.init = 16'h2222;
    LUT4 i13082_4_lut_4_lut (.A(n17289), .B(n26), .C(n30), .D(n25), 
         .Z(LOGIC_CLOCK_enable_69)) /* synthesis lut_function=((B (C (D)))+!A) */ ;
    defparam i13082_4_lut_4_lut.init = 16'hd555;
    LUT4 currPixel_7__bdd_4_lut (.A(currPixel[7]), .B(currPixel[0]), .C(currPixel[1]), 
         .D(n17392), .Z(n16803)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam currPixel_7__bdd_4_lut.init = 16'h0020;
    CCU2D add_107_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(currPWMCount[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n14003), .S1(currPWMCount_15__N_254[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_1.INIT0 = 16'hF000;
    defparam add_107_1.INIT1 = 16'h5555;
    defparam add_107_1.INJECT1_0 = "NO";
    defparam add_107_1.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_17 (.A0(currPWMCount_c[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14096), .S1(Matrix_CTRL_Out_c_2));
    defparam sub_989_add_2_17.INIT0 = 16'h5555;
    defparam sub_989_add_2_17.INIT1 = 16'h0000;
    defparam sub_989_add_2_17.INJECT1_0 = "NO";
    defparam sub_989_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_646 (.A(currPixel[7]), .B(n17289), .C(n15705), .D(n4_adj_2494), 
         .Z(PIXEL_CLOCK_enable_20)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(153[4] 189[11])
    defparam i1_4_lut_adj_646.init = 16'h5f5d;
    LUT4 i1_2_lut (.A(currPixel[1]), .B(currPixel[0]), .Z(n4_adj_2494)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(153[4] 189[11])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 currPixel_996_mux_6_i1_3_lut (.A(currPixel[0]), .B(n37[0]), .C(n1840), 
         .Z(n47[0])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_mux_6_i1_3_lut.init = 16'hc5c5;
    CCU2D sub_989_add_2_15 (.A0(currPWMCount_c[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount_c[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14095), .COUT(n14096));
    defparam sub_989_add_2_15.INIT0 = 16'h5555;
    defparam sub_989_add_2_15.INIT1 = 16'h5555;
    defparam sub_989_add_2_15.INJECT1_0 = "NO";
    defparam sub_989_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_13 (.A0(\currPWMCount[11] ), .B0(currPWMVal[11]), 
          .C0(GND_net), .D0(GND_net), .A1(\currPWMCount[12] ), .B1(currPWMVal[12]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14094), .COUT(n14095));
    defparam sub_989_add_2_13.INIT0 = 16'h5999;
    defparam sub_989_add_2_13.INIT1 = 16'h5999;
    defparam sub_989_add_2_13.INJECT1_0 = "NO";
    defparam sub_989_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_11 (.A0(currPWMCount[9]), .B0(currPWMVal[9]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[10]), .B1(currPWMVal[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14093), .COUT(n14094));
    defparam sub_989_add_2_11.INIT0 = 16'h5999;
    defparam sub_989_add_2_11.INIT1 = 16'h5999;
    defparam sub_989_add_2_11.INJECT1_0 = "NO";
    defparam sub_989_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_9 (.A0(currPWMCount[7]), .B0(currPWMVal[7]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[8]), .B1(currPWMVal[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14092), .COUT(n14093));
    defparam sub_989_add_2_9.INIT0 = 16'h5999;
    defparam sub_989_add_2_9.INIT1 = 16'h5999;
    defparam sub_989_add_2_9.INJECT1_0 = "NO";
    defparam sub_989_add_2_9.INJECT1_1 = "NO";
    CCU2D add_10507_15 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14257), .S1(BUS_VALID_N_110));
    defparam add_10507_15.INIT0 = 16'heeee;
    defparam add_10507_15.INIT1 = 16'h0000;
    defparam add_10507_15.INJECT1_0 = "NO";
    defparam add_10507_15.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_7 (.A0(\currPWMCount[5] ), .B0(currPWMVal[5]), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[6] ), .B1(currPWMVal[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14091), .COUT(n14092));
    defparam sub_989_add_2_7.INIT0 = 16'h5999;
    defparam sub_989_add_2_7.INIT1 = 16'h5999;
    defparam sub_989_add_2_7.INJECT1_0 = "NO";
    defparam sub_989_add_2_7.INJECT1_1 = "NO";
    CCU2D add_10507_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[18] ), .D0(lastAddress_31__N_1310), .A1(\BUS_currGrantID[0] ), 
          .B1(\BUS_currGrantID[1] ), .C1(GND_net), .D1(GND_net), .CIN(n14256), 
          .COUT(n14257));
    defparam add_10507_13.INIT0 = 16'hff20;
    defparam add_10507_13.INIT1 = 16'heeee;
    defparam add_10507_13.INJECT1_0 = "NO";
    defparam add_10507_13.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_5 (.A0(\currPWMCount[3] ), .B0(currPWMVal[3]), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[4] ), .B1(currPWMVal[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14090), .COUT(n14091));
    defparam sub_989_add_2_5.INIT0 = 16'h5999;
    defparam sub_989_add_2_5.INIT1 = 16'h5999;
    defparam sub_989_add_2_5.INJECT1_0 = "NO";
    defparam sub_989_add_2_5.INJECT1_1 = "NO";
    CCU2D add_10507_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[16] ), .D0(n18277), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[17] ), .D1(n18264), 
          .CIN(n14255), .COUT(n14256));
    defparam add_10507_11.INIT0 = 16'h00ce;
    defparam add_10507_11.INIT1 = 16'h00ce;
    defparam add_10507_11.INJECT1_0 = "NO";
    defparam add_10507_11.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_3 (.A0(\currPWMCount[1] ), .B0(currPWMVal[1]), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[2] ), .B1(currPWMVal[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14089), .COUT(n14090));
    defparam sub_989_add_2_3.INIT0 = 16'h5999;
    defparam sub_989_add_2_3.INIT1 = 16'h5999;
    defparam sub_989_add_2_3.INJECT1_0 = "NO";
    defparam sub_989_add_2_3.INJECT1_1 = "NO";
    CCU2D add_10507_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[14] ), .D0(n18262), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[15] ), .D1(n18271), 
          .CIN(n14254), .COUT(n14255));
    defparam add_10507_9.INIT0 = 16'h00ce;
    defparam add_10507_9.INIT1 = 16'h00ce;
    defparam add_10507_9.INJECT1_0 = "NO";
    defparam add_10507_9.INJECT1_1 = "NO";
    CCU2D sub_989_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(currPWMCount[0]), .B1(currPWMVal[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n14089));
    defparam sub_989_add_2_1.INIT0 = 16'h0000;
    defparam sub_989_add_2_1.INIT1 = 16'h5999;
    defparam sub_989_add_2_1.INJECT1_0 = "NO";
    defparam sub_989_add_2_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut_rep_281 (.A(n3296), .B(currPWMCount_c[13]), .C(currPWMCount_c[14]), 
         .D(currPWMCount_c[15]), .Z(n17289)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_rep_281.init = 16'hfffe;
    LUT4 currBit_3__I_0_164_i15_4_lut (.A(n15779), .B(n8_adj_2495), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_11)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(143[26:55])
    defparam currBit_3__I_0_164_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_164_i8_3_lut (.A(\BLUE[3] [8]), .B(\BLUE[3] [9]), 
         .C(currBit[0]), .Z(n8_adj_2495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(143[26:55])
    defparam currBit_3__I_0_164_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_165_i15_4_lut (.A(n15786), .B(n8_adj_2496), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_10)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(142[27:56])
    defparam currBit_3__I_0_165_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_165_i8_3_lut (.A(\GREEN[3] [8]), .B(\GREEN[3] [9]), 
         .C(currBit[0]), .Z(n8_adj_2496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(142[27:56])
    defparam currBit_3__I_0_165_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_166_i15_4_lut (.A(n15793), .B(n8_adj_2497), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_9)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(141[24:53])
    defparam currBit_3__I_0_166_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_166_i8_3_lut (.A(\RED[3] [8]), .B(\RED[3] [9]), 
         .C(currBit[0]), .Z(n8_adj_2497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(141[24:53])
    defparam currBit_3__I_0_166_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_167_i15_4_lut (.A(n15800), .B(n8_adj_2498), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_8)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(139[25:54])
    defparam currBit_3__I_0_167_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_167_i8_3_lut (.A(\BLUE[2] [8]), .B(\BLUE[2] [9]), 
         .C(currBit[0]), .Z(n8_adj_2498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(139[25:54])
    defparam currBit_3__I_0_167_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_168_i15_4_lut (.A(n15807), .B(n8_adj_2499), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_7)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(138[26:55])
    defparam currBit_3__I_0_168_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_168_i8_3_lut (.A(\GREEN[2] [8]), .B(\GREEN[2] [9]), 
         .C(currBit[0]), .Z(n8_adj_2499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(138[26:55])
    defparam currBit_3__I_0_168_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_169_i15_4_lut (.A(n15814), .B(n8_adj_2500), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_6)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(137[24:53])
    defparam currBit_3__I_0_169_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_169_i8_3_lut (.A(\RED[2] [8]), .B(\RED[2] [9]), 
         .C(currBit[0]), .Z(n8_adj_2500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(137[24:53])
    defparam currBit_3__I_0_169_i8_3_lut.init = 16'hcaca;
    FD1P3IX currPixel_996__i6 (.D(n37[6]), .SP(PIXEL_CLOCK_enable_20), .CD(n17365), 
            .CK(PIXEL_CLOCK), .Q(currPixel[6])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i6.GSR = "DISABLED";
    LUT4 currBit_3__I_0_170_i15_4_lut (.A(n15821), .B(n8_adj_2501), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_5)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(135[25:54])
    defparam currBit_3__I_0_170_i15_4_lut.init = 16'hca0a;
    FD1P3IX currPixel_996__i5 (.D(n37[5]), .SP(PIXEL_CLOCK_enable_20), .CD(n17365), 
            .CK(PIXEL_CLOCK), .Q(currPixel[5])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i5.GSR = "DISABLED";
    LUT4 currBit_3__I_0_170_i8_3_lut (.A(\BLUE[1] [8]), .B(\BLUE[1] [9]), 
         .C(currBit[0]), .Z(n8_adj_2501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(135[25:54])
    defparam currBit_3__I_0_170_i8_3_lut.init = 16'hcaca;
    CCU2D add_10507_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[12] ), .D0(n18272), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[13] ), .D1(n18266), 
          .CIN(n14253), .COUT(n14254));
    defparam add_10507_7.INIT0 = 16'h00ce;
    defparam add_10507_7.INIT1 = 16'h00ce;
    defparam add_10507_7.INJECT1_0 = "NO";
    defparam add_10507_7.INJECT1_1 = "NO";
    LUT4 currBit_3__I_0_171_i15_4_lut (.A(n15828), .B(n8_adj_2502), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_4)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(134[26:55])
    defparam currBit_3__I_0_171_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_171_i8_3_lut (.A(\GREEN[1] [8]), .B(\GREEN[1] [9]), 
         .C(currBit[0]), .Z(n8_adj_2502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(134[26:55])
    defparam currBit_3__I_0_171_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_172_i15_4_lut (.A(n15835), .B(n8_adj_2503), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_3)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(133[24:53])
    defparam currBit_3__I_0_172_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_172_i8_3_lut (.A(\RED[1] [8]), .B(\RED[1] [9]), 
         .C(currBit[0]), .Z(n8_adj_2503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(133[24:53])
    defparam currBit_3__I_0_172_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_173_i15_4_lut (.A(n15842), .B(n8_adj_2504), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_2)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(131[25:54])
    defparam currBit_3__I_0_173_i15_4_lut.init = 16'hca0a;
    CCU2D add_10507_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[10] ), .D0(n18269), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[11] ), .D1(n18273), 
          .CIN(n14252), .COUT(n14253));
    defparam add_10507_5.INIT0 = 16'hff31;
    defparam add_10507_5.INIT1 = 16'h00ce;
    defparam add_10507_5.INJECT1_0 = "NO";
    defparam add_10507_5.INJECT1_1 = "NO";
    LUT4 currBit_3__I_0_173_i8_3_lut (.A(\BLUE[0] [8]), .B(\BLUE[0] [9]), 
         .C(currBit[0]), .Z(n8_adj_2504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(131[25:54])
    defparam currBit_3__I_0_173_i8_3_lut.init = 16'hcaca;
    CCU2D add_10507_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[8] ), .D0(n18267), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[9] ), .D1(n18268), 
          .CIN(n14251), .COUT(n14252));
    defparam add_10507_3.INIT0 = 16'h00ce;
    defparam add_10507_3.INIT1 = 16'h00ce;
    defparam add_10507_3.INJECT1_0 = "NO";
    defparam add_10507_3.INJECT1_1 = "NO";
    CCU2D add_10507_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[7] ), 
          .D1(n18274), .COUT(n14251));
    defparam add_10507_1.INIT0 = 16'hF000;
    defparam add_10507_1.INIT1 = 16'h00ce;
    defparam add_10507_1.INJECT1_0 = "NO";
    defparam add_10507_1.INJECT1_1 = "NO";
    LUT4 currBit_3__I_0_174_i15_4_lut (.A(n15849), .B(n8_adj_2505), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_1)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(130[26:55])
    defparam currBit_3__I_0_174_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_174_i8_3_lut (.A(\GREEN[0] [8]), .B(\GREEN[0] [9]), 
         .C(currBit[0]), .Z(n8_adj_2505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(130[26:55])
    defparam currBit_3__I_0_174_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_184_i15_4_lut (.A(n15856), .B(n8_adj_2506), .C(currBit[3]), 
         .D(n17435), .Z(Matrix_DATA_Out_c_0)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(129[24:53])
    defparam currBit_3__I_0_184_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_184_i8_3_lut (.A(\RED[0] [8]), .B(\RED[0] [9]), 
         .C(currBit[0]), .Z(n8_adj_2506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(129[24:53])
    defparam currBit_3__I_0_184_i8_3_lut.init = 16'hcaca;
    LUT4 i12984_4_lut (.A(MATRIX_CURRROW[3]), .B(MATRIX_CURRROW[2]), .C(MATRIX_CURRROW[0]), 
         .D(n6_adj_2507), .Z(Matrix_LINE_SEL_Out_c_2)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(147[29:46])
    defparam i12984_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_adj_647 (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[4]), 
         .Z(n6_adj_2507)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(147[29:46])
    defparam i1_2_lut_adj_647.init = 16'heeee;
    LUT4 i6566_2_lut (.A(PIXEL_CLOCK), .B(MATRIX_CLKEN_LAT), .Z(Matrix_CTRL_Out_c_0)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(201[18:66])
    defparam i6566_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_307_3_lut (.A(currPixel[7]), .B(n17392), .C(currPixel[1]), 
         .Z(PIXEL_CLOCK_enable_5)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_307_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_648 (.A(currPixel[7]), .B(n17392), .C(currPixel[0]), 
         .D(currPixel[1]), .Z(PIXEL_CLOCK_enable_9)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_648.init = 16'h0200;
    LUT4 i2_2_lut_3_lut_4_lut (.A(currPixel[7]), .B(n17392), .C(currPixel[0]), 
         .D(currPixel[1]), .Z(PIXEL_CLOCK_enable_3)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3AX currPixel_996__i1 (.D(n47[1]), .SP(PIXEL_CLOCK_enable_20), .CK(PIXEL_CLOCK), 
            .Q(currPixel[1])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i1.GSR = "DISABLED";
    FD1S3AX currPixel_996__i7 (.D(n25_adj_2508), .CK(PIXEL_CLOCK), .Q(currPixel[7])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i7.GSR = "DISABLED";
    FD1P3IX currPixel_996__i4 (.D(n37[4]), .SP(PIXEL_CLOCK_enable_20), .CD(n17365), 
            .CK(PIXEL_CLOCK), .Q(currPixel[4])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i4.GSR = "DISABLED";
    PFUMX i10302 (.BLUT(n15474), .ALUT(n148), .C0(currBit[3]), .Z(n13454));
    LUT4 i1_2_lut_rep_345 (.A(currPixel[0]), .B(n17392), .Z(n17353)) /* synthesis lut_function=((B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i1_2_lut_rep_345.init = 16'hdddd;
    LUT4 i13057_2_lut_3_lut (.A(currPixel[0]), .B(n17392), .C(currPixel[1]), 
         .Z(MATRIX_ROWCLK_N_279)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i13057_2_lut_3_lut.init = 16'h0202;
    LUT4 i13108_2_lut_3_lut_4_lut (.A(currPixel[0]), .B(n17392), .C(currBit[0]), 
         .D(currPixel[1]), .Z(n10348)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i13108_2_lut_3_lut_4_lut.init = 16'h0200;
    FD1P3IX currPixel_996__i3 (.D(n37[3]), .SP(PIXEL_CLOCK_enable_20), .CD(n17365), 
            .CK(PIXEL_CLOCK), .Q(currPixel[3])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i3.GSR = "DISABLED";
    LUT4 i3843_2_lut_3_lut_4_lut (.A(currPixel[0]), .B(n17392), .C(currBit[3]), 
         .D(currPixel[1]), .Z(n7187)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i3843_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i12994_2_lut_rep_308_3_lut (.A(currPixel[0]), .B(n17392), .C(currPixel[1]), 
         .Z(PIXEL_CLOCK_N_293_enable_26)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i12994_2_lut_rep_308_3_lut.init = 16'h2020;
    LUT4 i3_2_lut_3_lut (.A(currPixel[0]), .B(n17392), .C(currPixel[7]), 
         .Z(PIXEL_CLOCK_enable_7)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i3_2_lut_3_lut.init = 16'h2020;
    LUT4 i3838_2_lut_3_lut_4_lut (.A(currPixel[0]), .B(n17392), .C(currBit[0]), 
         .D(currPixel[1]), .Z(n7190)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i3838_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i3839_2_lut_3_lut_4_lut (.A(currPixel[0]), .B(n17392), .C(currBit[2]), 
         .D(currPixel[1]), .Z(n7191)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(163[10:27])
    defparam i3839_2_lut_3_lut_4_lut.init = 16'h2000;
    L6MUX21 i12131 (.D0(n15791), .D1(n15792), .SD(currBit[2]), .Z(n15793));
    LUT4 i13078_2_lut_rep_346 (.A(currPixel[0]), .B(n17392), .Z(n17354)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(170[10:27])
    defparam i13078_2_lut_rep_346.init = 16'h1111;
    L6MUX21 i12138 (.D0(n15798), .D1(n15799), .SD(currBit[2]), .Z(n15800));
    LUT4 i2_3_lut_4_lut_adj_649 (.A(currPixel[0]), .B(n17392), .C(currPixel[7]), 
         .D(currPixel[1]), .Z(n14612)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(170[10:27])
    defparam i2_3_lut_4_lut_adj_649.init = 16'h0010;
    L6MUX21 i12145 (.D0(n15805), .D1(n15806), .SD(currBit[2]), .Z(n15807));
    L6MUX21 i12152 (.D0(n15812), .D1(n15813), .SD(currBit[2]), .Z(n15814));
    L6MUX21 i12159 (.D0(n15819), .D1(n15820), .SD(currBit[2]), .Z(n15821));
    L6MUX21 i12166 (.D0(n15826), .D1(n15827), .SD(currBit[2]), .Z(n15828));
    L6MUX21 i12173 (.D0(n15833), .D1(n15834), .SD(currBit[2]), .Z(n15835));
    FD1P3IX currPixel_996__i2 (.D(n37[2]), .SP(PIXEL_CLOCK_enable_20), .CD(n17365), 
            .CK(PIXEL_CLOCK), .Q(currPixel[2])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996__i2.GSR = "DISABLED";
    L6MUX21 i12180 (.D0(n15840), .D1(n15841), .SD(currBit[2]), .Z(n15842));
    L6MUX21 i12187 (.D0(n15847), .D1(n15848), .SD(currBit[2]), .Z(n15849));
    LUT4 n138_bdd_4_lut (.A(n138), .B(n139), .C(currBit[0]), .D(currBit[1]), 
         .Z(currPWMVal_15__N_205[10])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n138_bdd_4_lut.init = 16'h00ca;
    L6MUX21 i12194 (.D0(n15854), .D1(n15855), .SD(currBit[2]), .Z(n15856));
    L6MUX21 i12117 (.D0(n15777), .D1(n15778), .SD(currBit[2]), .Z(n15779));
    L6MUX21 i12124 (.D0(n15784), .D1(n15785), .SD(currBit[2]), .Z(n15786));
    CCU2D add_107_13 (.A0(\currPWMCount[11] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\currPWMCount[12] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14008), .COUT(n14009), .S0(currPWMCount_15__N_254[11]), 
          .S1(currPWMCount_15__N_254[12]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_13.INIT0 = 16'h5aaa;
    defparam add_107_13.INIT1 = 16'h5aaa;
    defparam add_107_13.INJECT1_0 = "NO";
    defparam add_107_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_454 (.A(currBit[2]), .B(currBit[3]), .Z(n17462)) /* synthesis lut_function=(!((B)+!A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_rep_454.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_3_lut (.A(currBit[2]), .B(currBit[3]), 
         .C(currBit[1]), .Z(currPWMCountMax_15__N_222[8])) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_3_lut_4_lut_4_lut_3_lut.init = 16'h2424;
    LUT4 i7_1_lut_rep_455 (.A(currPixel[1]), .Z(n17463)) /* synthesis lut_function=(!(A)) */ ;
    defparam i7_1_lut_rep_455.init = 16'h5555;
    LUT4 i1_4_lut_4_lut_adj_650 (.A(currPixel[1]), .B(n17289), .C(n15705), 
         .D(currPixel[0]), .Z(n15367)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_650.init = 16'h0f04;
    LUT4 i10330_3_lut_rep_456 (.A(\PWMArray[0] [12]), .B(\PWMArray[0] [10]), 
         .C(currBit[1]), .Z(n17464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10330_3_lut_rep_456.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(\PWMArray[0] [12]), .B(\PWMArray[0] [10]), .C(currBit[1]), 
         .D(currBit[3]), .Z(n4_c)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i1_2_lut_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_3_lut_adj_651 (.A(currBit[2]), .B(currBit[1]), .C(\PWMArray[0] [12]), 
         .Z(n15474)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_3_lut_adj_651.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_652 (.A(currBit[2]), .B(\PWMArray[0] [11]), 
         .C(currBit[3]), .Z(n139)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_3_lut_adj_652.init = 16'h4040;
    LUT4 i10339_4_lut_4_lut (.A(currBit[2]), .B(\PWMArray[0] [11]), .C(\PWMArray[0][9] ), 
         .D(currBit[1]), .Z(n13491)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10339_4_lut_4_lut.init = 16'h44a0;
    LUT4 i1_2_lut_rep_459 (.A(currBit[2]), .B(\PWMArray[0] [12]), .Z(n17467)) /* synthesis lut_function=(!(A+!(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_rep_459.init = 16'h4444;
    LUT4 i10337_4_lut_4_lut (.A(currBit[2]), .B(\PWMArray[0] [12]), .C(\PWMArray[0] [10]), 
         .D(currBit[1]), .Z(n13489)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10337_4_lut_4_lut.init = 16'h44a0;
    LUT4 VRAM_READ_ADDR_7__I_0_1_lut_rep_462 (.A(VRAM_READ_ADDR[7]), .Z(n17470)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(240[24:44])
    defparam VRAM_READ_ADDR_7__I_0_1_lut_rep_462.init = 16'h5555;
    CCU2D add_10510_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14209), 
          .S0(n2469));
    defparam add_10510_cout.INIT0 = 16'h0000;
    defparam add_10510_cout.INIT1 = 16'h0000;
    defparam add_10510_cout.INJECT1_0 = "NO";
    defparam add_10510_cout.INJECT1_1 = "NO";
    CCU2D add_10510_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14208), .COUT(n14209));
    defparam add_10510_21.INIT0 = 16'heeee;
    defparam add_10510_21.INIT1 = 16'heeee;
    defparam add_10510_21.INJECT1_0 = "NO";
    defparam add_10510_21.INJECT1_1 = "NO";
    CCU2D add_10510_19 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[17] ), .D0(n18264), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), .D1(lastAddress_31__N_1310), 
          .CIN(n14207), .COUT(n14208));
    defparam add_10510_19.INIT0 = 16'h00ce;
    defparam add_10510_19.INIT1 = 16'hff20;
    defparam add_10510_19.INJECT1_0 = "NO";
    defparam add_10510_19.INJECT1_1 = "NO";
    LUT4 i12191_3_lut (.A(\RED[0] [6]), .B(\RED[0] [7]), .C(currBit[0]), 
         .Z(n15853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12191_3_lut.init = 16'hcaca;
    CCU2D add_10510_17 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n18271), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16] ), .D1(n18277), 
          .CIN(n14206), .COUT(n14207));
    defparam add_10510_17.INIT0 = 16'h00ce;
    defparam add_10510_17.INIT1 = 16'h00ce;
    defparam add_10510_17.INJECT1_0 = "NO";
    defparam add_10510_17.INJECT1_1 = "NO";
    PFUMX i13412 (.BLUT(n17477), .ALUT(n17478), .C0(VRAM_READ_ADDR[7]), 
          .Z(VRAM_READ_ADDR_7__N_124));
    LUT4 i12190_3_lut (.A(\RED[0] [4]), .B(\RED[0] [5]), .C(currBit[0]), 
         .Z(n15852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12190_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_357 (.A(n15705), .B(currPixel[7]), .C(currPixel[1]), 
         .Z(n17365)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i2_3_lut_rep_357.init = 16'h4040;
    LUT4 i1_2_lut_4_lut_adj_653 (.A(n15705), .B(currPixel[7]), .C(currPixel[1]), 
         .D(currPixel[0]), .Z(n15359)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_4_lut_adj_653.init = 16'h4000;
    CCU2D add_10510_15 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n18266), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n18262), 
          .CIN(n14205), .COUT(n14206));
    defparam add_10510_15.INIT0 = 16'h00ce;
    defparam add_10510_15.INIT1 = 16'h00ce;
    defparam add_10510_15.INJECT1_0 = "NO";
    defparam add_10510_15.INJECT1_1 = "NO";
    LUT4 SpriteRead_yInSprite_7__N_597_7__I_0_i6_3_lut_3_lut_4_lut (.A(MATRIX_CURRROW[3]), 
         .B(n17408), .C(\SpriteRead_yValid_N_1158[2] ), .D(\SpriteRead_yValid_N_1158[3] ), 
         .Z(n6)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (B (C (D))+!B (C+(D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam SpriteRead_yInSprite_7__N_597_7__I_0_i6_3_lut_3_lut_4_lut.init = 16'hf990;
    LUT4 i1_2_lut_rep_291_3_lut_4_lut (.A(MATRIX_CURRROW[3]), .B(n17408), 
         .C(\SpriteRead_yValid_N_1158[4] ), .D(MATRIX_CURRROW[4]), .Z(n17299)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_rep_291_3_lut_4_lut.init = 16'h8778;
    LUT4 i12189_3_lut (.A(\RED[0] [2]), .B(\RED[0] [3]), .C(currBit[0]), 
         .Z(n15851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12189_3_lut.init = 16'hcaca;
    CCU2D add_10510_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n18273), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n18272), 
          .CIN(n14204), .COUT(n14205));
    defparam add_10510_13.INIT0 = 16'h00ce;
    defparam add_10510_13.INIT1 = 16'h00ce;
    defparam add_10510_13.INJECT1_0 = "NO";
    defparam add_10510_13.INJECT1_1 = "NO";
    LUT4 i12188_3_lut (.A(\RED[0] [0]), .B(\RED[0] [1]), .C(currBit[0]), 
         .Z(n15850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12188_3_lut.init = 16'hcaca;
    CCU2D add_10510_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[9] ), .D0(n18268), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n18269), 
          .CIN(n14203), .COUT(n14204));
    defparam add_10510_11.INIT0 = 16'h00ce;
    defparam add_10510_11.INIT1 = 16'hff31;
    defparam add_10510_11.INJECT1_0 = "NO";
    defparam add_10510_11.INJECT1_1 = "NO";
    CCU2D add_10510_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[7] ), .D0(n18274), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), .D1(n18267), 
          .CIN(n14202), .COUT(n14203));
    defparam add_10510_9.INIT0 = 16'hff31;
    defparam add_10510_9.INIT1 = 16'h00ce;
    defparam add_10510_9.INJECT1_0 = "NO";
    defparam add_10510_9.INJECT1_1 = "NO";
    CCU2D add_10510_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[5] ), .D0(n18265), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[6] ), .D1(n18276), 
          .CIN(n14201), .COUT(n14202));
    defparam add_10510_7.INIT0 = 16'h00ce;
    defparam add_10510_7.INIT1 = 16'h00ce;
    defparam add_10510_7.INJECT1_0 = "NO";
    defparam add_10510_7.INJECT1_1 = "NO";
    CCU2D add_10510_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[3] ), .D0(n17409), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[4] ), .D1(n18275), 
          .CIN(n14200), .COUT(n14201));
    defparam add_10510_5.INIT0 = 16'h00ce;
    defparam add_10510_5.INIT1 = 16'h00ce;
    defparam add_10510_5.INJECT1_0 = "NO";
    defparam add_10510_5.INJECT1_1 = "NO";
    CCU2D add_10510_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[1] ), .D0(n17423), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[2] ), .D1(n18263), 
          .CIN(n14199), .COUT(n14200));
    defparam add_10510_3.INIT0 = 16'h00ce;
    defparam add_10510_3.INIT1 = 16'h00ce;
    defparam add_10510_3.INJECT1_0 = "NO";
    defparam add_10510_3.INJECT1_1 = "NO";
    LUT4 i12184_3_lut (.A(\GREEN[0] [6]), .B(\GREEN[0] [7]), .C(currBit[0]), 
         .Z(n15846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12184_3_lut.init = 16'hcaca;
    LUT4 i12183_3_lut (.A(\GREEN[0] [4]), .B(\GREEN[0] [5]), .C(currBit[0]), 
         .Z(n15845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12183_3_lut.init = 16'hcaca;
    CCU2D add_10510_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[0] ), 
          .D1(n18261), .COUT(n14199));
    defparam add_10510_1.INIT0 = 16'hF000;
    defparam add_10510_1.INIT1 = 16'h00ce;
    defparam add_10510_1.INJECT1_0 = "NO";
    defparam add_10510_1.INJECT1_1 = "NO";
    LUT4 i12121_3_lut (.A(\GREEN[3] [6]), .B(\GREEN[3] [7]), .C(currBit[0]), 
         .Z(n15783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12121_3_lut.init = 16'hcaca;
    LUT4 i800_2_lut (.A(currBit[0]), .B(currBit[1]), .Z(n3)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(195[36:65])
    defparam i800_2_lut.init = 16'h6666;
    LUT4 i12177_3_lut (.A(\BLUE[0] [6]), .B(\BLUE[0] [7]), .C(currBit[0]), 
         .Z(n15839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12177_3_lut.init = 16'hcaca;
    LUT4 currPixel_996_mux_6_i2_3_lut (.A(currPixel[0]), .B(n37[1]), .C(n1840), 
         .Z(n47[1])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_996_mux_6_i2_3_lut.init = 16'hc5c5;
    LUT4 i13085_4_lut (.A(n15359), .B(n37[7]), .C(currPixel[7]), .D(n15367), 
         .Z(n25_adj_2508)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i13085_4_lut.init = 16'h4454;
    LUT4 i10309_4_lut_then_4_lut (.A(currBit[2]), .B(currBit[1]), .C(currBit[3]), 
         .D(\PWMArray[0][9] ), .Z(n17487)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10309_4_lut_then_4_lut.init = 16'h1808;
    LUT4 i10309_4_lut_else_4_lut (.A(currBit[2]), .B(currBit[1]), .C(currBit[3]), 
         .D(\PWMArray[0][9] ), .Z(n17486)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i10309_4_lut_else_4_lut.init = 16'h1000;
    LUT4 i1557_1_lut (.A(MATRIX_CURRROW[0]), .Z(\SpriteRead_yInSprite_7__N_597[0] )) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1557_1_lut.init = 16'h5555;
    LUT4 i2_3_lut_rep_296_4_lut (.A(n17329), .B(n17328), .C(n17458), .D(n15539), 
         .Z(n17304)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(275[55:66])
    defparam i2_3_lut_rep_296_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_adj_654 (.A(\PWMArray[0] [10]), .B(n13509), .Z(n161)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam i1_2_lut_adj_654.init = 16'h8888;
    LUT4 i3845_3_lut_4_lut (.A(n17353), .B(currPixel[1]), .C(currBit[3]), 
         .D(currBit[2]), .Z(n7196)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(183[10:27])
    defparam i3845_3_lut_4_lut.init = 16'h4440;
    LUT4 i1_2_lut_adj_655 (.A(\PWMArray[0] [11]), .B(n13509), .Z(n160)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam i1_2_lut_adj_655.init = 16'h8888;
    LUT4 i1_2_lut_adj_656 (.A(\PWMArray[0] [12]), .B(n13509), .Z(n159)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(281[3] 288[10])
    defparam i1_2_lut_adj_656.init = 16'h8888;
    LUT4 i1846_2_lut_4_lut (.A(n16803), .B(n17391), .C(currBit[3]), .D(MATRIX_CURRROW[0]), 
         .Z(n12[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(152[3] 190[10])
    defparam i1846_2_lut_4_lut.init = 16'h7f80;
    LUT4 i1_2_lut_then_4_lut (.A(currBit[1]), .B(currBit[3]), .C(currBit[2]), 
         .D(\PWMArray[0] [12]), .Z(n17493)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_then_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_rep_309_4_lut (.A(currBit[0]), .B(n17435), .C(currBit[3]), 
         .D(n16803), .Z(PIXEL_CLOCK_enable_13)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(66[9:16])
    defparam i2_3_lut_rep_309_4_lut.init = 16'hb000;
    LUT4 i5_4_lut_rep_384 (.A(n9), .B(n15633), .C(currPixel[7]), .D(currPixel[3]), 
         .Z(n17392)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(170[10:27])
    defparam i5_4_lut_rep_384.init = 16'hffef;
    LUT4 i1_2_lut_rep_343_4_lut (.A(n9), .B(n15633), .C(currPixel[7]), 
         .D(currPixel[3]), .Z(n17351)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(170[10:27])
    defparam i1_2_lut_rep_343_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_else_4_lut (.A(currBit[1]), .B(\PWMArray[0] [11]), .C(currBit[3]), 
         .D(currBit[2]), .Z(n17492)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_else_4_lut.init = 16'h0004;
    LUT4 i12119_3_lut (.A(\GREEN[3] [2]), .B(\GREEN[3] [3]), .C(currBit[0]), 
         .Z(n15781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12119_3_lut.init = 16'hcaca;
    LUT4 i12118_3_lut (.A(\GREEN[3] [0]), .B(\GREEN[3] [1]), .C(currBit[0]), 
         .Z(n15780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12118_3_lut.init = 16'hcaca;
    LUT4 i12126_3_lut (.A(\RED[3] [2]), .B(\RED[3] [3]), .C(currBit[0]), 
         .Z(n15788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12126_3_lut.init = 16'hcaca;
    PFUMX i12129 (.BLUT(n15787), .ALUT(n15788), .C0(currBit[1]), .Z(n15791));
    LUT4 i12176_3_lut (.A(\BLUE[0] [4]), .B(\BLUE[0] [5]), .C(currBit[0]), 
         .Z(n15838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12176_3_lut.init = 16'hcaca;
    LUT4 i12125_3_lut (.A(\RED[3] [0]), .B(\RED[3] [1]), .C(currBit[0]), 
         .Z(n15787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12125_3_lut.init = 16'hcaca;
    PFUMX i12130 (.BLUT(n15789), .ALUT(n15790), .C0(currBit[1]), .Z(n15792));
    LUT4 i12114_3_lut (.A(\BLUE[3] [6]), .B(\BLUE[3] [7]), .C(currBit[0]), 
         .Z(n15776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12114_3_lut.init = 16'hcaca;
    LUT4 i12113_3_lut (.A(\BLUE[3] [4]), .B(\BLUE[3] [5]), .C(currBit[0]), 
         .Z(n15775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12113_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_299_3_lut_4_lut (.A(MATRIX_CURRROW[2]), .B(n17452), 
         .C(\SpriteRead_yValid_N_1158[3] ), .D(MATRIX_CURRROW[3]), .Z(n17307)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1_2_lut_rep_299_3_lut_4_lut.init = 16'h8778;
    LUT4 i1580_2_lut_rep_318_3_lut_4_lut (.A(MATRIX_CURRROW[2]), .B(n17452), 
         .C(MATRIX_CURRROW[4]), .D(MATRIX_CURRROW[3]), .Z(n17326)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1580_2_lut_rep_318_3_lut_4_lut.init = 16'h78f0;
    PFUMX i12136 (.BLUT(n15794), .ALUT(n15795), .C0(currBit[1]), .Z(n15798));
    PFUMX i12137 (.BLUT(n15796), .ALUT(n15797), .C0(currBit[1]), .Z(n15799));
    PFUMX i12143 (.BLUT(n15801), .ALUT(n15802), .C0(currBit[1]), .Z(n15805));
    PFUMX i12144 (.BLUT(n15803), .ALUT(n15804), .C0(currBit[1]), .Z(n15806));
    PFUMX i12150 (.BLUT(n15808), .ALUT(n15809), .C0(currBit[1]), .Z(n15812));
    LUT4 i3_2_lut (.A(currPixel[5]), .B(currPixel[6]), .Z(n9)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(170[10:27])
    defparam i3_2_lut.init = 16'heeee;
    PFUMX i12151 (.BLUT(n15810), .ALUT(n15811), .C0(currBit[1]), .Z(n15813));
    PFUMX i12157 (.BLUT(n15815), .ALUT(n15816), .C0(currBit[1]), .Z(n15819));
    LUT4 i12112_3_lut (.A(\BLUE[3] [2]), .B(\BLUE[3] [3]), .C(currBit[0]), 
         .Z(n15774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12112_3_lut.init = 16'hcaca;
    PFUMX i12158 (.BLUT(n15817), .ALUT(n15818), .C0(currBit[1]), .Z(n15820));
    LUT4 i12111_3_lut (.A(\BLUE[3] [0]), .B(\BLUE[3] [1]), .C(currBit[0]), 
         .Z(n15773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12111_3_lut.init = 16'hcaca;
    PFUMX i12164 (.BLUT(n15822), .ALUT(n15823), .C0(currBit[1]), .Z(n15826));
    LUT4 i12182_3_lut (.A(\GREEN[0] [2]), .B(\GREEN[0] [3]), .C(currBit[0]), 
         .Z(n15844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12182_3_lut.init = 16'hcaca;
    LUT4 i12181_3_lut (.A(\GREEN[0] [0]), .B(\GREEN[0] [1]), .C(currBit[0]), 
         .Z(n15843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12181_3_lut.init = 16'hcaca;
    PFUMX i12165 (.BLUT(n15824), .ALUT(n15825), .C0(currBit[1]), .Z(n15827));
    PFUMX i12171 (.BLUT(n15829), .ALUT(n15830), .C0(currBit[1]), .Z(n15833));
    PFUMX i12172 (.BLUT(n15831), .ALUT(n15832), .C0(currBit[1]), .Z(n15834));
    PFUMX i12178 (.BLUT(n15836), .ALUT(n15837), .C0(currBit[1]), .Z(n15840));
    PFUMX i12179 (.BLUT(n15838), .ALUT(n15839), .C0(currBit[1]), .Z(n15841));
    Outputbuffer VRam (.VRAM_DATA({VRAM_DATA}), .GND_net(GND_net), .n17470(n17470), 
            .\VRAM_ADDR[8] (\VRAM_ADDR[8] ), .\VRAM_ADDR[7] (\VRAM_ADDR[7] ), 
            .\VRAM_ADDR[6] (\VRAM_ADDR[6] ), .\VRAM_ADDR[5] (\VRAM_ADDR[5] ), 
            .\VRAM_ADDR[4] (\VRAM_ADDR[4] ), .\VRAM_ADDR[3] (\VRAM_ADDR[3] ), 
            .\VRAM_ADDR[2] (\VRAM_ADDR[2] ), .\VRAM_ADDR[1] (\VRAM_ADDR[1] ), 
            .\VRAM_ADDR[0] (\VRAM_ADDR[0] ), .\VRAM_READ_ADDR[7] (VRAM_READ_ADDR[7]), 
            .\currPixel[6] (currPixel[6]), .\currPixel[5] (currPixel[5]), 
            .\currPixel[4] (currPixel[4]), .\currPixel[3] (currPixel[3]), 
            .\currPixel[2] (currPixel[2]), .\currPixel[1] (currPixel[1]), 
            .\currPixel[0] (currPixel[0]), .VRAM_WC(VRAM_WC), .PIXEL_CLOCK_N_293(PIXEL_CLOCK_N_293), 
            .VCC_net(VCC_net), .VRAM_WE(VRAM_WE), .VRAM_DATA_OUT({VRAM_DATA_OUT}), 
            .\BLUE[3] ({\BLUE[3] }), .\BLUE[2] ({\BLUE[2] }), .\BLUE[1] ({\BLUE[1] }), 
            .\BLUE[0] ({\BLUE[0] }), .\RED[3] ({\RED[3] }), .\RED[2] ({\RED[2] }), 
            .\RED[1] ({\RED[1] }), .\RED[0] ({\RED[0] }), .\GREEN[3] ({\GREEN[3] }), 
            .\GREEN[2] ({\GREEN[2] }), .\GREEN[1] ({\GREEN[1] }), .\GREEN[0] ({\GREEN[0] })) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    
endmodule
//
// Verilog Description of module Outputbuffer
//

module Outputbuffer (VRAM_DATA, GND_net, n17470, \VRAM_ADDR[8] , \VRAM_ADDR[7] , 
            \VRAM_ADDR[6] , \VRAM_ADDR[5] , \VRAM_ADDR[4] , \VRAM_ADDR[3] , 
            \VRAM_ADDR[2] , \VRAM_ADDR[1] , \VRAM_ADDR[0] , \VRAM_READ_ADDR[7] , 
            \currPixel[6] , \currPixel[5] , \currPixel[4] , \currPixel[3] , 
            \currPixel[2] , \currPixel[1] , \currPixel[0] , VRAM_WC, 
            PIXEL_CLOCK_N_293, VCC_net, VRAM_WE, VRAM_DATA_OUT, \BLUE[3] , 
            \BLUE[2] , \BLUE[1] , \BLUE[0] , \RED[3] , \RED[2] , \RED[1] , 
            \RED[0] , \GREEN[3] , \GREEN[2] , \GREEN[1] , \GREEN[0] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [29:0]VRAM_DATA;
    input GND_net;
    input n17470;
    input \VRAM_ADDR[8] ;
    input \VRAM_ADDR[7] ;
    input \VRAM_ADDR[6] ;
    input \VRAM_ADDR[5] ;
    input \VRAM_ADDR[4] ;
    input \VRAM_ADDR[3] ;
    input \VRAM_ADDR[2] ;
    input \VRAM_ADDR[1] ;
    input \VRAM_ADDR[0] ;
    input \VRAM_READ_ADDR[7] ;
    input \currPixel[6] ;
    input \currPixel[5] ;
    input \currPixel[4] ;
    input \currPixel[3] ;
    input \currPixel[2] ;
    input \currPixel[1] ;
    input \currPixel[0] ;
    input VRAM_WC;
    input PIXEL_CLOCK_N_293;
    input VCC_net;
    input VRAM_WE;
    output [29:0]VRAM_DATA_OUT;
    output [9:0]\BLUE[3] ;
    output [9:0]\BLUE[2] ;
    output [9:0]\BLUE[1] ;
    output [9:0]\BLUE[0] ;
    output [9:0]\RED[3] ;
    output [9:0]\RED[2] ;
    output [9:0]\RED[1] ;
    output [9:0]\RED[0] ;
    output [9:0]\GREEN[3] ;
    output [9:0]\GREEN[2] ;
    output [9:0]\GREEN[1] ;
    output [9:0]\GREEN[0] ;
    
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(91[8:15])
    wire PIXEL_CLOCK_N_293 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(88[9:22])
    
    DP8KC Outputbuffer_0_14_0 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[28]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[29]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[28]), .DOA1(VRAM_DATA_OUT[29]), 
          .DOB0(\BLUE[0] [8]), .DOB1(\BLUE[0] [9]), .DOB2(\BLUE[1] [8]), 
          .DOB3(\BLUE[1] [9]), .DOB4(\BLUE[2] [8]), .DOB5(\BLUE[2] [9]), 
          .DOB6(\BLUE[3] [8]), .DOB7(\BLUE[3] [9])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_14_0.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_14_0.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_14_0.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_14_0.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_14_0.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_14_0.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_14_0.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_14_0.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_14_0.GSR = "ENABLED";
    defparam Outputbuffer_0_14_0.RESETMODE = "SYNC";
    defparam Outputbuffer_0_14_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_14_0.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_14_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_14_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_1_13 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[2]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[3]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[2]), .DOA1(VRAM_DATA_OUT[3]), 
          .DOB0(\RED[0] [2]), .DOB1(\RED[0] [3]), .DOB2(\RED[1] [2]), 
          .DOB3(\RED[1] [3]), .DOB4(\RED[2] [2]), .DOB5(\RED[2] [3]), 
          .DOB6(\RED[3] [2]), .DOB7(\RED[3] [3])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_1_13.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_1_13.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_1_13.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_1_13.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_1_13.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_1_13.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_1_13.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_1_13.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_1_13.GSR = "ENABLED";
    defparam Outputbuffer_0_1_13.RESETMODE = "SYNC";
    defparam Outputbuffer_0_1_13.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_1_13.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_1_13.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_1_13.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_0_14 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[0]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[1]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[0]), .DOA1(VRAM_DATA_OUT[1]), 
          .DOB0(\RED[0] [0]), .DOB1(\RED[0] [1]), .DOB2(\RED[1] [0]), 
          .DOB3(\RED[1] [1]), .DOB4(\RED[2] [0]), .DOB5(\RED[2] [1]), 
          .DOB6(\RED[3] [0]), .DOB7(\RED[3] [1])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_0_14.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_0_14.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_0_14.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_0_14.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_0_14.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_0_14.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_0_14.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_0_14.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_0_14.GSR = "ENABLED";
    defparam Outputbuffer_0_0_14.RESETMODE = "SYNC";
    defparam Outputbuffer_0_0_14.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_0_14.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_0_14.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_0_14.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_2_12 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[4]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[5]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[4]), .DOA1(VRAM_DATA_OUT[5]), 
          .DOB0(\RED[0] [4]), .DOB1(\RED[0] [5]), .DOB2(\RED[1] [4]), 
          .DOB3(\RED[1] [5]), .DOB4(\RED[2] [4]), .DOB5(\RED[2] [5]), 
          .DOB6(\RED[3] [4]), .DOB7(\RED[3] [5])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_2_12.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_2_12.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_2_12.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_2_12.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_2_12.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_2_12.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_2_12.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_2_12.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_2_12.GSR = "ENABLED";
    defparam Outputbuffer_0_2_12.RESETMODE = "SYNC";
    defparam Outputbuffer_0_2_12.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_2_12.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_2_12.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_2_12.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_3_11 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[6]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[7]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[6]), .DOA1(VRAM_DATA_OUT[7]), 
          .DOB0(\RED[0] [6]), .DOB1(\RED[0] [7]), .DOB2(\RED[1] [6]), 
          .DOB3(\RED[1] [7]), .DOB4(\RED[2] [6]), .DOB5(\RED[2] [7]), 
          .DOB6(\RED[3] [6]), .DOB7(\RED[3] [7])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_3_11.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_3_11.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_3_11.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_3_11.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_3_11.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_3_11.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_3_11.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_3_11.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_3_11.GSR = "ENABLED";
    defparam Outputbuffer_0_3_11.RESETMODE = "SYNC";
    defparam Outputbuffer_0_3_11.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_3_11.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_3_11.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_3_11.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_4_10 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[8]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[9]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[8]), .DOA1(VRAM_DATA_OUT[9]), 
          .DOB0(\RED[0] [8]), .DOB1(\RED[0] [9]), .DOB2(\RED[1] [8]), 
          .DOB3(\RED[1] [9]), .DOB4(\RED[2] [8]), .DOB5(\RED[2] [9]), 
          .DOB6(\RED[3] [8]), .DOB7(\RED[3] [9])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_4_10.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_4_10.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_4_10.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_4_10.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_4_10.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_4_10.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_4_10.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_4_10.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_4_10.GSR = "ENABLED";
    defparam Outputbuffer_0_4_10.RESETMODE = "SYNC";
    defparam Outputbuffer_0_4_10.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_4_10.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_4_10.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_4_10.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_5_9 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[10]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[11]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[10]), .DOA1(VRAM_DATA_OUT[11]), 
          .DOB0(\GREEN[0] [0]), .DOB1(\GREEN[0] [1]), .DOB2(\GREEN[1] [0]), 
          .DOB3(\GREEN[1] [1]), .DOB4(\GREEN[2] [0]), .DOB5(\GREEN[2] [1]), 
          .DOB6(\GREEN[3] [0]), .DOB7(\GREEN[3] [1])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_5_9.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_5_9.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_5_9.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_5_9.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_5_9.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_5_9.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_5_9.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_5_9.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_5_9.GSR = "ENABLED";
    defparam Outputbuffer_0_5_9.RESETMODE = "SYNC";
    defparam Outputbuffer_0_5_9.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_5_9.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_5_9.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_5_9.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_6_8 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[12]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[13]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[12]), .DOA1(VRAM_DATA_OUT[13]), 
          .DOB0(\GREEN[0] [2]), .DOB1(\GREEN[0] [3]), .DOB2(\GREEN[1] [2]), 
          .DOB3(\GREEN[1] [3]), .DOB4(\GREEN[2] [2]), .DOB5(\GREEN[2] [3]), 
          .DOB6(\GREEN[3] [2]), .DOB7(\GREEN[3] [3])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_6_8.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_6_8.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_6_8.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_6_8.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_6_8.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_6_8.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_6_8.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_6_8.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_6_8.GSR = "ENABLED";
    defparam Outputbuffer_0_6_8.RESETMODE = "SYNC";
    defparam Outputbuffer_0_6_8.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_6_8.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_6_8.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_6_8.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_7_7 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[14]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[15]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[14]), .DOA1(VRAM_DATA_OUT[15]), 
          .DOB0(\GREEN[0] [4]), .DOB1(\GREEN[0] [5]), .DOB2(\GREEN[1] [4]), 
          .DOB3(\GREEN[1] [5]), .DOB4(\GREEN[2] [4]), .DOB5(\GREEN[2] [5]), 
          .DOB6(\GREEN[3] [4]), .DOB7(\GREEN[3] [5])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_7_7.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_7_7.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_7_7.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_7_7.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_7_7.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_7_7.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_7_7.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_7_7.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_7_7.GSR = "ENABLED";
    defparam Outputbuffer_0_7_7.RESETMODE = "SYNC";
    defparam Outputbuffer_0_7_7.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_7_7.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_7_7.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_7_7.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_8_6 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[16]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[17]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[16]), .DOA1(VRAM_DATA_OUT[17]), 
          .DOB0(\GREEN[0] [6]), .DOB1(\GREEN[0] [7]), .DOB2(\GREEN[1] [6]), 
          .DOB3(\GREEN[1] [7]), .DOB4(\GREEN[2] [6]), .DOB5(\GREEN[2] [7]), 
          .DOB6(\GREEN[3] [6]), .DOB7(\GREEN[3] [7])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_8_6.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_8_6.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_8_6.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_8_6.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_8_6.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_8_6.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_8_6.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_8_6.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_8_6.GSR = "ENABLED";
    defparam Outputbuffer_0_8_6.RESETMODE = "SYNC";
    defparam Outputbuffer_0_8_6.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_8_6.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_8_6.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_8_6.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_9_5 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[18]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[19]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[18]), .DOA1(VRAM_DATA_OUT[19]), 
          .DOB0(\GREEN[0] [8]), .DOB1(\GREEN[0] [9]), .DOB2(\GREEN[1] [8]), 
          .DOB3(\GREEN[1] [9]), .DOB4(\GREEN[2] [8]), .DOB5(\GREEN[2] [9]), 
          .DOB6(\GREEN[3] [8]), .DOB7(\GREEN[3] [9])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_9_5.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_9_5.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_9_5.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_9_5.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_9_5.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_9_5.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_9_5.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_9_5.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_9_5.GSR = "ENABLED";
    defparam Outputbuffer_0_9_5.RESETMODE = "SYNC";
    defparam Outputbuffer_0_9_5.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_9_5.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_9_5.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_9_5.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_10_4 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[20]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[21]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[20]), .DOA1(VRAM_DATA_OUT[21]), 
          .DOB0(\BLUE[0] [0]), .DOB1(\BLUE[0] [1]), .DOB2(\BLUE[1] [0]), 
          .DOB3(\BLUE[1] [1]), .DOB4(\BLUE[2] [0]), .DOB5(\BLUE[2] [1]), 
          .DOB6(\BLUE[3] [0]), .DOB7(\BLUE[3] [1])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_10_4.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_10_4.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_10_4.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_10_4.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_10_4.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_10_4.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_10_4.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_10_4.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_10_4.GSR = "ENABLED";
    defparam Outputbuffer_0_10_4.RESETMODE = "SYNC";
    defparam Outputbuffer_0_10_4.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_10_4.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_10_4.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_10_4.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_11_3 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[22]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[23]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[22]), .DOA1(VRAM_DATA_OUT[23]), 
          .DOB0(\BLUE[0] [2]), .DOB1(\BLUE[0] [3]), .DOB2(\BLUE[1] [2]), 
          .DOB3(\BLUE[1] [3]), .DOB4(\BLUE[2] [2]), .DOB5(\BLUE[2] [3]), 
          .DOB6(\BLUE[3] [2]), .DOB7(\BLUE[3] [3])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_11_3.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_11_3.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_11_3.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_11_3.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_11_3.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_11_3.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_11_3.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_11_3.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_11_3.GSR = "ENABLED";
    defparam Outputbuffer_0_11_3.RESETMODE = "SYNC";
    defparam Outputbuffer_0_11_3.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_11_3.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_11_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_11_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_12_2 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[24]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[25]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[24]), .DOA1(VRAM_DATA_OUT[25]), 
          .DOB0(\BLUE[0] [4]), .DOB1(\BLUE[0] [5]), .DOB2(\BLUE[1] [4]), 
          .DOB3(\BLUE[1] [5]), .DOB4(\BLUE[2] [4]), .DOB5(\BLUE[2] [5]), 
          .DOB6(\BLUE[3] [4]), .DOB7(\BLUE[3] [5])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_12_2.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_12_2.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_12_2.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_12_2.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_12_2.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_12_2.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_12_2.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_12_2.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_12_2.GSR = "ENABLED";
    defparam Outputbuffer_0_12_2.RESETMODE = "SYNC";
    defparam Outputbuffer_0_12_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_12_2.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_12_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_12_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC Outputbuffer_0_13_1 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(VRAM_DATA[26]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(VRAM_DATA[27]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(\VRAM_ADDR[0] ), 
          .ADA2(\VRAM_ADDR[1] ), .ADA3(\VRAM_ADDR[2] ), .ADA4(\VRAM_ADDR[3] ), 
          .ADA5(\VRAM_ADDR[4] ), .ADA6(\VRAM_ADDR[5] ), .ADA7(\VRAM_ADDR[6] ), 
          .ADA8(\VRAM_ADDR[7] ), .ADA9(\VRAM_ADDR[8] ), .ADA10(n17470), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(VRAM_WC), .WEA(VRAM_WE), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(\currPixel[0] ), .ADB4(\currPixel[1] ), 
          .ADB5(\currPixel[2] ), .ADB6(\currPixel[3] ), .ADB7(\currPixel[4] ), 
          .ADB8(\currPixel[5] ), .ADB9(\currPixel[6] ), .ADB10(\VRAM_READ_ADDR[7] ), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(PIXEL_CLOCK_N_293), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(VRAM_DATA_OUT[26]), .DOA1(VRAM_DATA_OUT[27]), 
          .DOB0(\BLUE[0] [6]), .DOB1(\BLUE[0] [7]), .DOB2(\BLUE[1] [6]), 
          .DOB3(\BLUE[1] [7]), .DOB4(\BLUE[2] [6]), .DOB5(\BLUE[2] [7]), 
          .DOB6(\BLUE[3] [6]), .DOB7(\BLUE[3] [7])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=250, LSE_RLINE=250 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(250[8:20])
    defparam Outputbuffer_0_13_1.DATA_WIDTH_A = 2;
    defparam Outputbuffer_0_13_1.DATA_WIDTH_B = 9;
    defparam Outputbuffer_0_13_1.REGMODE_A = "OUTREG";
    defparam Outputbuffer_0_13_1.REGMODE_B = "OUTREG";
    defparam Outputbuffer_0_13_1.CSDECODE_A = "0b000";
    defparam Outputbuffer_0_13_1.CSDECODE_B = "0b000";
    defparam Outputbuffer_0_13_1.WRITEMODE_A = "NORMAL";
    defparam Outputbuffer_0_13_1.WRITEMODE_B = "NORMAL";
    defparam Outputbuffer_0_13_1.GSR = "ENABLED";
    defparam Outputbuffer_0_13_1.RESETMODE = "SYNC";
    defparam Outputbuffer_0_13_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_13_1.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_13_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Outputbuffer_0_13_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PLL
//

module PLL (LOGIC_CLOCK_N_57, LOGIC_CLOCK, CLK_c, PIXEL_CLOCK, GND_net, 
            PIXEL_CLOCK_N_293) /* synthesis NGD_DRC_MASK=1 */ ;
    output LOGIC_CLOCK_N_57;
    output LOGIC_CLOCK;
    input CLK_c;
    output PIXEL_CLOCK;
    input GND_net;
    output PIXEL_CLOCK_N_293;
    
    wire LOGIC_CLOCK_N_57 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire CLK_c /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    wire PIXEL_CLOCK /* synthesis SET_AS_NETWORK=PIXEL_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(43[8:19])
    wire PIXEL_CLOCK_N_293 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(88[9:22])
    
    INV i13875 (.A(LOGIC_CLOCK), .Z(LOGIC_CLOCK_N_57));
    EHXPLLJ PLLInst_0 (.CLKI(CLK_c), .CLKFB(LOGIC_CLOCK), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(LOGIC_CLOCK), .CLKOS(PIXEL_CLOCK)) /* synthesis FREQUENCY_PIN_CLKOS="35.416667", FREQUENCY_PIN_CLKOP="141.666667", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="8", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=244, LSE_RLINE=244 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(244[10:13])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 17;
    defparam PLLInst_0.CLKOP_DIV = 4;
    defparam PLLInst_0.CLKOS_DIV = 16;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 3;
    defparam PLLInst_0.CLKOS_CPHASE = 15;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    INV i13876 (.A(PIXEL_CLOCK), .Z(PIXEL_CLOCK_N_293));
    
endmodule
//
// Verilog Description of module MatrixBusHandler
//

module MatrixBusHandler (VRAM_DATA_OUT, GND_net, LOGIC_CLOCK, n17458, 
            n17411, n18270, n17382, lastAddress_31__N_1338, \BUS_DATA_INTERNAL[7] , 
            yOffset, n17339, n17333, n17332, n17331, BUS_data, n4305, 
            n4306, n4307, n4308, \state[0] , \BUS_DATA_INTERNAL[6] , 
            n17276, n17314, n17334, n17321, n17312, \BUS_DATA_INTERNAL[5] , 
            \SpriteRead_yInSprite_7__N_597[0] , \VRAM_ADDR[0] , \BUS_DATA_INTERNAL[4] , 
            n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, 
            n4616, n4617, n4618, n4619, n4573, n4574, n4575, n4576, 
            n4591, n17381, lastAddress_31__N_1323, n4577, n4578, n4579, 
            n4580, n4581, n4582, n4583, n4584, n4592, n4593, n4594, 
            n4595, n4625, n4596, n4597, n4598, n4599, n4600, n4601, 
            n4602, n4603, n2877, \BUS_DATA_INTERNAL[3] , n4557, n4558, 
            n4559, n4560, n4590, n4561, n4562, n4563, n4564, n17373, 
            lastAddress_31__N_1413, n2878, \BUS_DATA_INTERNAL[2] , n2879, 
            \BUS_DATA_INTERNAL[1] , SpriteRead_yValid_N_1158, n2880, \BUS_DATA_INTERNAL[0] , 
            n4604, n4605, n4606, n4607, VRAM_WC, n8, VRAM_DATA, 
            \BUS_ADDR_INTERNAL[0] , n4355, n4356, n4357, n4358, n4460, 
            n4461, n4462, n4463, n4565, n4566, n4567, n4568, Sprite_pointers_N_1123, 
            VCC_net, n4250, n4251, n4252, n4253, n17342, n17310, 
            n4569, n4570, n4571, n4572, n4585, n4586, n4587, n4588, 
            n4620, n4621, n4622, n4623, n4503, n4504, n4505, n4506, 
            \Sprite_readData2[10] , n4507, n4508, n4509, n4510, n17371, 
            lastAddress_31__N_1337, \Sprite_readData2[11] , \Sprite_readData2[12] , 
            \Sprite_readData2[13] , n4511, n4512, n4513, n4514, n4468, 
            n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, 
            n4477, n4478, n4479, n18280, \Sprite_readData2[14] , \Sprite_readData2[15] , 
            latchMode, n17343, n4487, n4488, n4489, n4490, xOffset, 
            VRAM_WE, \state[1] , n4491, n4492, n4493, n4494, n4495, 
            n4496, n4497, n4498, n4452, n4453, n4454, n4455, n17366, 
            MATRIX_CURRROW, \BUS_ADDR_INTERNAL[3] , \BUS_currGrantID[0] , 
            \BUS_currGrantID[1] , \BUS_ADDR_INTERNAL[3]_adj_2 , n17453, 
            n17326, \BUS_ADDR_INTERNAL[14] , \BUS_ADDR_INTERNAL[14]_adj_3 , 
            n17383, \BUS_ADDR_INTERNAL[2] , \BUS_ADDR_INTERNAL[2]_adj_4 , 
            \BUS_ADDR_INTERNAL[17] , \BUS_ADDR_INTERNAL[17]_adj_5 , n18260, 
            n17272, \BUS_ADDR_INTERNAL[5] , \BUS_ADDR_INTERNAL[5]_adj_6 , 
            n17380, n4456, n4457, n4458, n4459, \BUS_ADDR_INTERNAL[13] , 
            \BUS_ADDR_INTERNAL[13]_adj_7 , n17379, \BUS_ADDR_INTERNAL[8] , 
            \BUS_ADDR_INTERNAL[8]_adj_8 , n17378, \BUS_ADDR_INTERNAL[9] , 
            \BUS_ADDR_INTERNAL[9]_adj_9 , n17376, \BUS_ADDR_INTERNAL[4] , 
            \BUS_ADDR_INTERNAL[4]_adj_10 , n17375, n17275, \state[1]_adj_11 , 
            n17434, n17457, n15469, \BUS_ADDR_INTERNAL[6] , \BUS_ADDR_INTERNAL[6]_adj_12 , 
            n17374, \BUS_ADDR_INTERNAL[7] , \BUS_ADDR_INTERNAL[7]_adj_13 , 
            \BUS_ADDR_INTERNAL[12] , \BUS_ADDR_INTERNAL[12]_adj_14 , n17377, 
            n17407, \BUS_ADDR_INTERNAL[16] , \BUS_ADDR_INTERNAL[16]_adj_15 , 
            n17362, \BUS_ADDR_INTERNAL[15] , \BUS_ADDR_INTERNAL[15]_adj_16 , 
            n17355, \state[3] , \yOffset[3] , \yOffset[2] , \yOffset[1] , 
            n16084, n16085, n4499, n4500, n4501, n4502, n16097, 
            n16098, n16107, n16108, n33, \BUS_ADDR_INTERNAL[0]_adj_17 , 
            n17385, n16114, n16115, n4464, n4465, n4466, n4467, 
            n4480, n4481, n4482, n4483, n4515, n4516, n4517, n4518, 
            n9891, n4398, n4399, n4400, n4401, BUS_DONE_OUT_N_1051, 
            n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, 
            n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
            n4371, n4372, n4373, n4374, n4382, n4383, n4384, n4385, 
            n4386, n4387, n4388, n4389, n16121, n16122, n4390, 
            n4391, n4392, n4393, n4347, n4348, n4349, n4350, n4351, 
            n4352, n4353, n4354, n16126, n16127, n16128, n16129, 
            n16130, n16131, n4394, n4395, n4396, n4397, n16132, 
            n16133, n4359, n4360, n4361, n4362, n4375, n4376, 
            n4377, n4378, n17329, n17327, n16141, n16142, n4410, 
            n4411, n4412, n4413, n4293, n4294, n4295, n4296, n4297, 
            n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4258, 
            n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
            n4267, n4268, n4269, n4277, n4278, n4279, n4280, n4281, 
            n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4242, 
            n4243, n4244, n4245, n4246, n4247, n4248, n4249, n17279, 
            n17274, n16143, n16144, n4289, n4290, n4291, n4292, 
            n16145, n16146, n4254, n4255, n4256, n4257, n4270, 
            n4271, n4272, n4273, n16147, n16148, n16156, n16157, 
            Sprite_pointers_N_1136, n17287, n16158, n16159, SpriteRead_yInSprite, 
            LOGIC_CLOCK_enable_52, \SpriteRead_yValid_N_1158[1] , n16160, 
            n16161, n16162, n16163, n16171, n16172, n18264, \BUS_ADDR_INTERNAL[18] , 
            lastAddress_31__N_1310, n18271, n18277, n18266, n18262, 
            n16173, n16174, n16175, n16176, \BUS_ADDR_INTERNAL[11] , 
            n18273, n18272, n16177, n16178, n18268, \BUS_ADDR_INTERNAL[10] , 
            n18269, n18267, n15749, n15750, n16186, n16187, n16188, 
            n16189, n16190, n16191, \BUS_currGrantID_3__N_74[0] , n17408, 
            n17368, n16192, n16193, n17452, n16201, n16202, n16203, 
            n16204, n16205, n16206, n16207, n16208, \BUS_ADDR_INTERNAL[18]_derived_1 , 
            n2504, n15752, n15753, lastAddress_31__N_1425, n17384, 
            n6250, n17311, n15755, n15756, n15758, n15759, n15761, 
            n15762, n16216, n16217, n16218, n16219, n16220, n16221, 
            n16222, n16223, reset, state_7__N_345, \Sprite_readAddr_13__N_752[13] , 
            n17313, \Sprite_readAddr_13__N_752[11] , \Sprite_readAddr_13__N_752[12] , 
            \Sprite_readAddr_13__N_752[9] , \Sprite_readAddr_13__N_752[10] , 
            n15764, n15765, n16231, n16232, n16234, n16235, \Sprite_readAddr_13__N_752[7] , 
            \Sprite_readAddr_13__N_752[8] , \Sprite_readAddr_13__N_752[5] , 
            \Sprite_readAddr_13__N_752[6] , \Sprite_readAddr_13__N_752[3] , 
            \Sprite_readAddr_13__N_752[4] , \Sprite_readAddr_13__N_752[1] , 
            \Sprite_readAddr_13__N_752[2] , n16237, n16238, \Sprite_readAddr_13__N_752[0] , 
            n17256, n16240, n16241, n16243, n16244, n16246, n16247, 
            n16251, n16252, n16256, n16257, n16259, n16260, n16262, 
            n16263, n15767, n15768, n16265, n16266, n15770, n15771, 
            n16270, n16271, n16275, n16276, n16278, n16279, n16281, 
            n16282, \VRAM_ADDR[1] , \VRAM_ADDR[2] , \VRAM_ADDR[3] , 
            \VRAM_ADDR[4] , \VRAM_ADDR[5] , \VRAM_ADDR[6] , \VRAM_ADDR[7] , 
            \VRAM_ADDR[8] , \BUS_ADDR_INTERNAL[1] , \BUS_ADDR_INTERNAL[10]_adj_18 , 
            \BUS_ADDR_INTERNAL[11]_adj_19 , n16284, n16285, n16287, 
            n16288, n17337, n17325, \BUS_addr[10] , \BUS_addr[11] , 
            n17335, n17338, \xOffset[2] , \xOffset[3] , n9, n16290, 
            n16291, n17340, n15655, n16293, n16294, n15436, n2642, 
            n16298, n16299, n16303, n16304, n16306, n16307, n16309, 
            n16310, n16312, n16313, n16315, n16316, n16320, n16321, 
            n4, n17305, n17298, n63, n63_adj_20, n16325, n16326, 
            n16328, n16329, n16331, n16332, n16334, n16335, n16337, 
            n16338, lastAddress_31__N_1434, n17302, n17309, n17308, 
            n16340, n16341, \currSprite_size[6] , \currSprite_size[7] , 
            lastAddress_31__N_1401, \currSprite_size[4] , \currSprite_size[5] , 
            lastAddress_31__N_1336, n17304, n7, n18276, n18274, \currSprite_size[2] , 
            \currSprite_size[3] , n18275, n18265, n18263, n17409, 
            n17423, n18259, n17394, \currSprite_size[1] , lastAddress_31__N_1422, 
            \MDM_data[8] , \otherData[9] , n15539, n17328, n6340, 
            SRAM_WE_N_1254, \lastAddress[18] , n46, lastAddress_31__N_1431, 
            lastAddress_31__N_1383, lastAddress_31__N_1325, lastAddress_31__N_1334, 
            lastAddress_31__N_1326, lastAddress_31__N_1404, lastAddress_31__N_1333, 
            lastAddress_31__N_1335, lastAddress_31__N_1330, lastAddress_31__N_1419, 
            lastAddress_31__N_1407, lastAddress_31__N_1395, lastAddress_31__N_1386, 
            lastAddress_31__N_1331, lastAddress_31__N_1389, lastAddress_31__N_1398, 
            lastAddress_31__N_1328, lastAddress_31__N_1392, lastAddress_31__N_1327, 
            lastAddress_31__N_1428, lastAddress_31__N_1339, lastAddress_31__N_1332, 
            lastAddress_31__N_1329, lastAddress_31__N_1324, lastAddress_31__N_1340, 
            lastAddress_31__N_1416, lastAddress_31__N_1410, n14584, \SpriteRead_yValid_N_1158[4] , 
            n17299, n17307, n15549, \SpriteRead_yValid_N_1158[0] , n15571, 
            n8_adj_21, WRITE_DONE, n10346, n17456, n17344, RED_WRITE, 
            GREEN_WRITE, LOGIC_CLOCK_N_57, n17387, BLUE_WRITE, ALPHA_WRITE);
    input [29:0]VRAM_DATA_OUT;
    input GND_net;
    input LOGIC_CLOCK;
    input n17458;
    input n17411;
    input n18270;
    output n17382;
    output lastAddress_31__N_1338;
    output \BUS_DATA_INTERNAL[7] ;
    output [7:0]yOffset;
    input n17339;
    output n17333;
    input n17332;
    input n17331;
    input [15:0]BUS_data;
    output n4305;
    output n4306;
    output n4307;
    output n4308;
    output \state[0] ;
    output \BUS_DATA_INTERNAL[6] ;
    output n17276;
    input n17314;
    input n17334;
    input n17321;
    input n17312;
    output \BUS_DATA_INTERNAL[5] ;
    input \SpriteRead_yInSprite_7__N_597[0] ;
    output \VRAM_ADDR[0] ;
    output \BUS_DATA_INTERNAL[4] ;
    output n4608;
    output n4609;
    output n4610;
    output n4611;
    output n4612;
    output n4613;
    output n4614;
    output n4615;
    output n4616;
    output n4617;
    output n4618;
    output n4619;
    output n4573;
    output n4574;
    output n4575;
    output n4576;
    input n4591;
    output n17381;
    output lastAddress_31__N_1323;
    output n4577;
    output n4578;
    output n4579;
    output n4580;
    output n4581;
    output n4582;
    output n4583;
    output n4584;
    output n4592;
    output n4593;
    output n4594;
    output n4595;
    input n4625;
    output n4596;
    output n4597;
    output n4598;
    output n4599;
    output n4600;
    output n4601;
    output n4602;
    output n4603;
    input n2877;
    output \BUS_DATA_INTERNAL[3] ;
    output n4557;
    output n4558;
    output n4559;
    output n4560;
    input n4590;
    output n4561;
    output n4562;
    output n4563;
    output n4564;
    output n17373;
    output lastAddress_31__N_1413;
    input n2878;
    output \BUS_DATA_INTERNAL[2] ;
    input n2879;
    output \BUS_DATA_INTERNAL[1] ;
    output [7:0]SpriteRead_yValid_N_1158;
    input n2880;
    output \BUS_DATA_INTERNAL[0] ;
    output n4604;
    output n4605;
    output n4606;
    output n4607;
    output VRAM_WC;
    input n8;
    output [29:0]VRAM_DATA;
    output \BUS_ADDR_INTERNAL[0] ;
    output n4355;
    output n4356;
    output n4357;
    output n4358;
    output n4460;
    output n4461;
    output n4462;
    output n4463;
    output n4565;
    output n4566;
    output n4567;
    output n4568;
    output Sprite_pointers_N_1123;
    input VCC_net;
    output n4250;
    output n4251;
    output n4252;
    output n4253;
    input n17342;
    input n17310;
    output n4569;
    output n4570;
    output n4571;
    output n4572;
    output n4585;
    output n4586;
    output n4587;
    output n4588;
    output n4620;
    output n4621;
    output n4622;
    output n4623;
    output n4503;
    output n4504;
    output n4505;
    output n4506;
    output \Sprite_readData2[10] ;
    output n4507;
    output n4508;
    output n4509;
    output n4510;
    output n17371;
    output lastAddress_31__N_1337;
    output \Sprite_readData2[11] ;
    output \Sprite_readData2[12] ;
    output \Sprite_readData2[13] ;
    output n4511;
    output n4512;
    output n4513;
    output n4514;
    output n4468;
    output n4469;
    output n4470;
    output n4471;
    output n4472;
    output n4473;
    output n4474;
    output n4475;
    output n4476;
    output n4477;
    output n4478;
    output n4479;
    input n18280;
    output \Sprite_readData2[14] ;
    output \Sprite_readData2[15] ;
    output [3:0]latchMode;
    input n17343;
    output n4487;
    output n4488;
    output n4489;
    output n4490;
    output [7:0]xOffset;
    output VRAM_WE;
    output \state[1] ;
    output n4491;
    output n4492;
    output n4493;
    output n4494;
    output n4495;
    output n4496;
    output n4497;
    output n4498;
    output n4452;
    output n4453;
    output n4454;
    output n4455;
    input n17366;
    input [4:0]MATRIX_CURRROW;
    input \BUS_ADDR_INTERNAL[3] ;
    input \BUS_currGrantID[0] ;
    input \BUS_currGrantID[1] ;
    output \BUS_ADDR_INTERNAL[3]_adj_2 ;
    input n17453;
    input n17326;
    output \BUS_ADDR_INTERNAL[14] ;
    input \BUS_ADDR_INTERNAL[14]_adj_3 ;
    output n17383;
    output \BUS_ADDR_INTERNAL[2] ;
    input \BUS_ADDR_INTERNAL[2]_adj_4 ;
    output \BUS_ADDR_INTERNAL[17] ;
    input \BUS_ADDR_INTERNAL[17]_adj_5 ;
    input n18260;
    output n17272;
    output \BUS_ADDR_INTERNAL[5] ;
    input \BUS_ADDR_INTERNAL[5]_adj_6 ;
    output n17380;
    output n4456;
    output n4457;
    output n4458;
    output n4459;
    output \BUS_ADDR_INTERNAL[13] ;
    input \BUS_ADDR_INTERNAL[13]_adj_7 ;
    output n17379;
    output \BUS_ADDR_INTERNAL[8] ;
    input \BUS_ADDR_INTERNAL[8]_adj_8 ;
    output n17378;
    output \BUS_ADDR_INTERNAL[9] ;
    input \BUS_ADDR_INTERNAL[9]_adj_9 ;
    output n17376;
    output \BUS_ADDR_INTERNAL[4] ;
    input \BUS_ADDR_INTERNAL[4]_adj_10 ;
    output n17375;
    output n17275;
    input \state[1]_adj_11 ;
    input n17434;
    input n17457;
    output n15469;
    output \BUS_ADDR_INTERNAL[6] ;
    input \BUS_ADDR_INTERNAL[6]_adj_12 ;
    output n17374;
    output \BUS_ADDR_INTERNAL[7] ;
    input \BUS_ADDR_INTERNAL[7]_adj_13 ;
    output \BUS_ADDR_INTERNAL[12] ;
    input \BUS_ADDR_INTERNAL[12]_adj_14 ;
    output n17377;
    input n17407;
    output \BUS_ADDR_INTERNAL[16] ;
    input \BUS_ADDR_INTERNAL[16]_adj_15 ;
    output n17362;
    output \BUS_ADDR_INTERNAL[15] ;
    input \BUS_ADDR_INTERNAL[15]_adj_16 ;
    output n17355;
    output \state[3] ;
    output \yOffset[3] ;
    output \yOffset[2] ;
    output \yOffset[1] ;
    input n16084;
    input n16085;
    output n4499;
    output n4500;
    output n4501;
    output n4502;
    input n16097;
    input n16098;
    input n16107;
    input n16108;
    input n33;
    input \BUS_ADDR_INTERNAL[0]_adj_17 ;
    output n17385;
    input n16114;
    input n16115;
    output n4464;
    output n4465;
    output n4466;
    output n4467;
    output n4480;
    output n4481;
    output n4482;
    output n4483;
    output n4515;
    output n4516;
    output n4517;
    output n4518;
    input n9891;
    output n4398;
    output n4399;
    output n4400;
    output n4401;
    input BUS_DONE_OUT_N_1051;
    output n4402;
    output n4403;
    output n4404;
    output n4405;
    output n4406;
    output n4407;
    output n4408;
    output n4409;
    output n4363;
    output n4364;
    output n4365;
    output n4366;
    output n4367;
    output n4368;
    output n4369;
    output n4370;
    output n4371;
    output n4372;
    output n4373;
    output n4374;
    output n4382;
    output n4383;
    output n4384;
    output n4385;
    output n4386;
    output n4387;
    output n4388;
    output n4389;
    input n16121;
    input n16122;
    output n4390;
    output n4391;
    output n4392;
    output n4393;
    output n4347;
    output n4348;
    output n4349;
    output n4350;
    output n4351;
    output n4352;
    output n4353;
    output n4354;
    input n16126;
    input n16127;
    input n16128;
    input n16129;
    input n16130;
    input n16131;
    output n4394;
    output n4395;
    output n4396;
    output n4397;
    input n16132;
    input n16133;
    output n4359;
    output n4360;
    output n4361;
    output n4362;
    output n4375;
    output n4376;
    output n4377;
    output n4378;
    output n17329;
    input n17327;
    input n16141;
    input n16142;
    output n4410;
    output n4411;
    output n4412;
    output n4413;
    output n4293;
    output n4294;
    output n4295;
    output n4296;
    output n4297;
    output n4298;
    output n4299;
    output n4300;
    output n4301;
    output n4302;
    output n4303;
    output n4304;
    output n4258;
    output n4259;
    output n4260;
    output n4261;
    output n4262;
    output n4263;
    output n4264;
    output n4265;
    output n4266;
    output n4267;
    output n4268;
    output n4269;
    output n4277;
    output n4278;
    output n4279;
    output n4280;
    output n4281;
    output n4282;
    output n4283;
    output n4284;
    output n4285;
    output n4286;
    output n4287;
    output n4288;
    output n4242;
    output n4243;
    output n4244;
    output n4245;
    output n4246;
    output n4247;
    output n4248;
    output n4249;
    input n17279;
    output n17274;
    input n16143;
    input n16144;
    output n4289;
    output n4290;
    output n4291;
    output n4292;
    input n16145;
    input n16146;
    output n4254;
    output n4255;
    output n4256;
    output n4257;
    output n4270;
    output n4271;
    output n4272;
    output n4273;
    input n16147;
    input n16148;
    input n16156;
    input n16157;
    input Sprite_pointers_N_1136;
    output n17287;
    input n16158;
    input n16159;
    output [7:0]SpriteRead_yInSprite;
    input LOGIC_CLOCK_enable_52;
    output \SpriteRead_yValid_N_1158[1] ;
    input n16160;
    input n16161;
    input n16162;
    input n16163;
    input n16171;
    input n16172;
    input n18264;
    input \BUS_ADDR_INTERNAL[18] ;
    input lastAddress_31__N_1310;
    input n18271;
    input n18277;
    input n18266;
    input n18262;
    input n16173;
    input n16174;
    input n16175;
    input n16176;
    input \BUS_ADDR_INTERNAL[11] ;
    input n18273;
    input n18272;
    input n16177;
    input n16178;
    input n18268;
    input \BUS_ADDR_INTERNAL[10] ;
    input n18269;
    input n18267;
    input n15749;
    input n15750;
    input n16186;
    input n16187;
    input n16188;
    input n16189;
    input n16190;
    input n16191;
    output \BUS_currGrantID_3__N_74[0] ;
    input n17408;
    input n17368;
    input n16192;
    input n16193;
    input n17452;
    input n16201;
    input n16202;
    input n16203;
    input n16204;
    input n16205;
    input n16206;
    input n16207;
    input n16208;
    input \BUS_ADDR_INTERNAL[18]_derived_1 ;
    output n2504;
    input n15752;
    input n15753;
    output lastAddress_31__N_1425;
    input n17384;
    input n6250;
    output n17311;
    input n15755;
    input n15756;
    input n15758;
    input n15759;
    input n15761;
    input n15762;
    input n16216;
    input n16217;
    input n16218;
    input n16219;
    input n16220;
    input n16221;
    input n16222;
    input n16223;
    output reset;
    output state_7__N_345;
    input \Sprite_readAddr_13__N_752[13] ;
    input n17313;
    input \Sprite_readAddr_13__N_752[11] ;
    input \Sprite_readAddr_13__N_752[12] ;
    input \Sprite_readAddr_13__N_752[9] ;
    input \Sprite_readAddr_13__N_752[10] ;
    input n15764;
    input n15765;
    input n16231;
    input n16232;
    input n16234;
    input n16235;
    input \Sprite_readAddr_13__N_752[7] ;
    input \Sprite_readAddr_13__N_752[8] ;
    input \Sprite_readAddr_13__N_752[5] ;
    input \Sprite_readAddr_13__N_752[6] ;
    input \Sprite_readAddr_13__N_752[3] ;
    input \Sprite_readAddr_13__N_752[4] ;
    input \Sprite_readAddr_13__N_752[1] ;
    input \Sprite_readAddr_13__N_752[2] ;
    input n16237;
    input n16238;
    input \Sprite_readAddr_13__N_752[0] ;
    input n17256;
    input n16240;
    input n16241;
    input n16243;
    input n16244;
    input n16246;
    input n16247;
    input n16251;
    input n16252;
    input n16256;
    input n16257;
    input n16259;
    input n16260;
    input n16262;
    input n16263;
    input n15767;
    input n15768;
    input n16265;
    input n16266;
    input n15770;
    input n15771;
    input n16270;
    input n16271;
    input n16275;
    input n16276;
    input n16278;
    input n16279;
    input n16281;
    input n16282;
    output \VRAM_ADDR[1] ;
    output \VRAM_ADDR[2] ;
    output \VRAM_ADDR[3] ;
    output \VRAM_ADDR[4] ;
    output \VRAM_ADDR[5] ;
    output \VRAM_ADDR[6] ;
    output \VRAM_ADDR[7] ;
    output \VRAM_ADDR[8] ;
    output \BUS_ADDR_INTERNAL[1] ;
    output \BUS_ADDR_INTERNAL[10]_adj_18 ;
    output \BUS_ADDR_INTERNAL[11]_adj_19 ;
    input n16284;
    input n16285;
    input n16287;
    input n16288;
    input n17337;
    input n17325;
    input \BUS_addr[10] ;
    input \BUS_addr[11] ;
    input n17335;
    input n17338;
    output \xOffset[2] ;
    output \xOffset[3] ;
    output n9;
    input n16290;
    input n16291;
    input n17340;
    input n15655;
    input n16293;
    input n16294;
    input n15436;
    output n2642;
    input n16298;
    input n16299;
    input n16303;
    input n16304;
    input n16306;
    input n16307;
    input n16309;
    input n16310;
    input n16312;
    input n16313;
    input n16315;
    input n16316;
    input n16320;
    input n16321;
    input n4;
    input n17305;
    input n17298;
    input n63;
    input n63_adj_20;
    input n16325;
    input n16326;
    input n16328;
    input n16329;
    input n16331;
    input n16332;
    input n16334;
    input n16335;
    input n16337;
    input n16338;
    output lastAddress_31__N_1434;
    input n17302;
    input n17309;
    input n17308;
    input n16340;
    input n16341;
    output \currSprite_size[6] ;
    output \currSprite_size[7] ;
    output lastAddress_31__N_1401;
    output \currSprite_size[4] ;
    output \currSprite_size[5] ;
    output lastAddress_31__N_1336;
    input n17304;
    output n7;
    input n18276;
    input n18274;
    output \currSprite_size[2] ;
    output \currSprite_size[3] ;
    input n18275;
    input n18265;
    input n18263;
    input n17409;
    input n17423;
    input n18259;
    output n17394;
    output \currSprite_size[1] ;
    output lastAddress_31__N_1422;
    output \MDM_data[8] ;
    output \otherData[9] ;
    output n15539;
    output n17328;
    output n6340;
    input SRAM_WE_N_1254;
    input \lastAddress[18] ;
    output n46;
    output lastAddress_31__N_1431;
    output lastAddress_31__N_1383;
    output lastAddress_31__N_1325;
    output lastAddress_31__N_1334;
    output lastAddress_31__N_1326;
    output lastAddress_31__N_1404;
    output lastAddress_31__N_1333;
    output lastAddress_31__N_1335;
    output lastAddress_31__N_1330;
    output lastAddress_31__N_1419;
    output lastAddress_31__N_1407;
    output lastAddress_31__N_1395;
    output lastAddress_31__N_1386;
    output lastAddress_31__N_1331;
    output lastAddress_31__N_1389;
    output lastAddress_31__N_1398;
    output lastAddress_31__N_1328;
    output lastAddress_31__N_1392;
    output lastAddress_31__N_1327;
    output lastAddress_31__N_1428;
    output lastAddress_31__N_1339;
    output lastAddress_31__N_1332;
    output lastAddress_31__N_1329;
    output lastAddress_31__N_1324;
    output lastAddress_31__N_1340;
    output lastAddress_31__N_1416;
    output lastAddress_31__N_1410;
    output n14584;
    output \SpriteRead_yValid_N_1158[4] ;
    input n17299;
    input n17307;
    input n15549;
    output \SpriteRead_yValid_N_1158[0] ;
    input n15571;
    input n8_adj_21;
    input WRITE_DONE;
    input n10346;
    input n17456;
    input n17344;
    output [8:0]RED_WRITE;
    output [8:0]GREEN_WRITE;
    input LOGIC_CLOCK_N_57;
    input n17387;
    output [8:0]BLUE_WRITE;
    output [8:0]ALPHA_WRITE;
    
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire lastReadRow_2_derived_5 /* synthesis is_clock=1, SET_AS_NETWORK=\MDM/lastReadRow[2]_derived_5 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(89[9:20])
    wire offsetLatchClockOrd /* synthesis is_clock=1, SET_AS_NETWORK=\MDM/offsetLatchClockOrd */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(93[9:28])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(91[8:15])
    wire Sprite_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[9:23])
    wire SpriteLut_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(203[9:26])
    wire SpriteLut_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(202[9:27])
    wire GR_WR_CLK /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(162[9:18])
    wire Sprite_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(179[9:24])
    wire LOGIC_CLOCK_N_57 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    wire [9:0]RED_OUT_9__N_768;
    
    wire mfco, mult_10u_9u_0_pp_0_10, mult_10u_9u_0_pp_0_9, mco_3, mult_10u_9u_0_pp_0_8, 
        mult_10u_9u_0_pp_0_7, mco_2, n14063;
    wire [9:0]currAddress_17__N_742;
    wire [31:0]currAddress;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(108[9:20])
    
    wire n14064, mult_10u_9u_0_pp_0_6, mult_10u_9u_0_pp_0_5, mco_1;
    wire [7:0]currSprite;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(190[9:19])
    
    wire LOGIC_CLOCK_enable_88;
    wire [7:0]n37;
    
    wire co_mult_9u_9u_0_1_4, co_mult_9u_9u_0_1_5, s_mult_9u_9u_0_1_13, 
        s_mult_9u_9u_0_1_14, mult_9u_9u_0_pp_2_14, mult_9u_9u_0_pp_2_13, 
        mult_9u_9u_0_pp_3_14, mult_9u_9u_0_pp_3_13, mult_10u_9u_0_pp_0_4, 
        mult_10u_9u_0_pp_0_3, mco;
    wire [18:0]GREEN_OUT_9__N_650;
    
    wire mult_10u_9u_0_pp_0_2, mult_10u_9u_0_cin_lr_0, co_t_mult_10u_9u_0_3_5, 
        mult_10u_9u_0_pp_4_17, s_mult_10u_9u_0_2_17, s_mult_10u_9u_0_2_18, 
        n59, n62;
    wire [7:0]state;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(87[9:14])
    
    wire n95, co_mult_9u_9u_0_1_3, s_mult_9u_9u_0_1_11, s_mult_9u_9u_0_1_12, 
        mult_9u_9u_0_pp_2_12, mult_9u_9u_0_pp_2_11, mult_9u_9u_0_pp_3_12, 
        mult_9u_9u_0_pp_3_11, co_mult_9u_9u_0_1_2, s_mult_9u_9u_0_1_9, 
        s_mult_9u_9u_0_1_10, mult_9u_9u_0_pp_2_10, mult_9u_9u_0_pp_2_9, 
        mult_9u_9u_0_pp_3_10, mult_9u_9u_0_pp_3_9, co_mult_9u_9u_0_1_1, 
        s_mult_9u_9u_0_1_7, s_mult_9u_9u_0_1_8, mult_9u_9u_0_pp_2_8, mult_9u_9u_0_pp_2_7, 
        mult_9u_9u_0_pp_3_8, mult_9u_9u_0_pp_3_7, co_t_mult_10u_9u_0_3_4, 
        mult_10u_9u_0_pp_4_15, mult_10u_9u_0_pp_4_16, s_mult_10u_9u_0_2_15, 
        s_mult_10u_9u_0_2_16, mult_9u_9u_0_pp_3_6, s_mult_9u_9u_0_1_6, 
        mult_9u_9u_0_pp_2_6, co_mult_9u_9u_0_0_6, s_mult_9u_9u_0_0_13, 
        co_t_mult_10u_9u_0_3_3, mult_10u_9u_0_pp_4_13, mult_10u_9u_0_pp_4_14, 
        s_mult_10u_9u_0_2_13, s_mult_10u_9u_0_2_14, co_t_mult_10u_9u_0_3_2, 
        mult_10u_9u_0_pp_4_11, mult_10u_9u_0_pp_4_12, s_mult_10u_9u_0_2_11, 
        s_mult_10u_9u_0_2_12, co_mult_9u_9u_0_0_5, s_mult_9u_9u_0_0_11, 
        s_mult_9u_9u_0_0_12, mult_9u_9u_0_pp_1_12, mult_9u_9u_0_pp_1_11, 
        co_t_mult_10u_9u_0_3_1, mult_10u_9u_0_pp_4_9, mult_10u_9u_0_pp_4_10, 
        s_mult_10u_9u_0_2_9, s_mult_10u_9u_0_2_10, mult_10u_9u_0_pp_4_8, 
        s_mult_10u_9u_0_2_8, co_mult_9u_9u_0_0_4, s_mult_9u_9u_0_0_9, 
        s_mult_9u_9u_0_0_10, mult_9u_9u_0_pp_0_10, mult_9u_9u_0_pp_0_9, 
        mult_9u_9u_0_pp_1_10, mult_9u_9u_0_pp_1_9, co_mult_10u_9u_0_2_7, 
        s_mult_10u_9u_0_1_17, s_mult_10u_9u_0_1_18, co_mult_10u_9u_0_2_6, 
        s_mult_10u_9u_0_1_15, s_mult_10u_9u_0_1_16, s_mult_10u_9u_0_0_15, 
        co_mult_10u_9u_0_2_5, s_mult_10u_9u_0_1_13, s_mult_10u_9u_0_1_14, 
        s_mult_10u_9u_0_0_13, s_mult_10u_9u_0_0_14, co_mult_10u_9u_0_2_4, 
        s_mult_10u_9u_0_1_11, s_mult_10u_9u_0_1_12, s_mult_10u_9u_0_0_11, 
        s_mult_10u_9u_0_0_12, co_mult_10u_9u_0_2_3, s_mult_10u_9u_0_1_9, 
        s_mult_10u_9u_0_1_10, s_mult_10u_9u_0_0_9, s_mult_10u_9u_0_0_10, 
        co_mult_10u_9u_0_2_2, s_mult_10u_9u_0_1_7, s_mult_10u_9u_0_1_8, 
        s_mult_10u_9u_0_0_7, s_mult_10u_9u_0_0_8, co_mult_10u_9u_0_2_1, 
        s_mult_10u_9u_0_1_6, s_mult_10u_9u_0_0_5, s_mult_10u_9u_0_0_6, 
        mult_10u_9u_0_pp_2_5, LOGIC_CLOCK_enable_33, LOGIC_CLOCK_enable_113, 
        mult_10u_9u_0_pp_2_4, s_mult_10u_9u_0_0_4, co_mult_10u_9u_0_1_6, 
        mult_10u_9u_0_pp_3_17, co_mult_9u_9u_0_0_3, s_mult_9u_9u_0_0_7, 
        s_mult_9u_9u_0_0_8, mult_9u_9u_0_pp_0_8, mult_9u_9u_0_pp_0_7, 
        mult_9u_9u_0_pp_1_8, mult_9u_9u_0_pp_1_7;
    wire [15:0]GR_WR_DOUT_16;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(158[9:22])
    
    wire LOGIC_CLOCK_enable_79;
    wire [9:0]GR_WR_DOUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(157[9:19])
    wire [17:0]RED_OUT_9__N_632;
    
    wire co_t_mult_9u_9u_0_3_1, mult_9u_9u_0_pp_4_9, mult_9u_9u_0_pp_4_10, 
        s_mult_9u_9u_0_2_9, s_mult_9u_9u_0_2_10, co_t_mult_9u_9u_0_3_2, 
        co_mult_9u_9u_0_0_2, s_mult_9u_9u_0_0_5, s_mult_9u_9u_0_0_6, mult_9u_9u_0_pp_0_6, 
        mult_9u_9u_0_pp_0_5, mult_9u_9u_0_pp_1_6, mult_9u_9u_0_pp_1_5, 
        co_mult_10u_9u_0_1_5, mult_10u_9u_0_pp_2_15, mult_10u_9u_0_pp_3_16, 
        mult_10u_9u_0_pp_3_15, co_mult_10u_9u_0_1_4, mult_10u_9u_0_pp_2_14, 
        mult_10u_9u_0_pp_2_13, mult_10u_9u_0_pp_3_14, mult_10u_9u_0_pp_3_13;
    wire [15:0]otherData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(121[9:18])
    wire [7:0]n2872;
    
    wire n1985;
    wire [7:0]yOffset_pre;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(95[9:20])
    
    wire n4040, n4041, n4042, n4043, n4380, n4311;
    wire [8:0]RED_READ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(209[9:17])
    wire [8:0]ALPHA_READ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(212[9:19])
    
    wire mult_9u_9u_0_pp_4_8, s_mult_9u_9u_0_2_8, co_mult_10u_9u_0_1_3, 
        mult_10u_9u_0_pp_2_12, mult_10u_9u_0_pp_2_11, mult_10u_9u_0_pp_3_12, 
        mult_10u_9u_0_pp_3_11;
    wire [7:0]state_7__N_336;
    wire [8:0]GREEN_READ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(210[9:19])
    
    wire mult_9u_9u_0_pp_4_8_adj_1880, mult_10u_9u_0_pp_4_8_adj_1881;
    wire [8:0]BLUE_READ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(211[9:18])
    
    wire mult_9u_9u_0_pp_4_8_adj_1882, co_mult_10u_9u_0_1_2, mult_10u_9u_0_pp_2_10, 
        mult_10u_9u_0_pp_2_9, mult_10u_9u_0_pp_3_10, mult_10u_9u_0_pp_3_9, 
        latchForce, LOGIC_CLOCK_enable_4, co_mult_10u_9u_0_1_1, mult_10u_9u_0_pp_2_8, 
        mult_10u_9u_0_pp_2_7, mult_10u_9u_0_pp_3_8, mult_10u_9u_0_pp_3_7, 
        co_mult_9u_9u_0_0_1, s_mult_9u_9u_0_0_4, mult_9u_9u_0_pp_0_4, 
        mult_9u_9u_0_pp_0_3, mult_9u_9u_0_pp_1_4, mult_9u_9u_0_pp_1_3, 
        mult_10u_9u_0_pp_3_6, mult_10u_9u_0_pp_2_6, co_mult_10u_9u_0_0_7, 
        co_mult_10u_9u_0_0_6, mult_10u_9u_0_pp_1_13;
    wire [7:0]currValue;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(110[9:18])
    wire [15:0]otherData2;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(175[9:19])
    
    wire co_mult_10u_9u_0_0_5, mult_10u_9u_0_pp_0_11, mult_10u_9u_0_pp_1_12, 
        mult_10u_9u_0_pp_1_11, mult_9u_9u_0_pp_1_2, mult_9u_9u_0_pp_0_2;
    wire [3:0]currColor;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(107[9:18])
    
    wire n7210;
    wire [3:0]n3;
    
    wire n17273, n4415;
    wire [4:0]lastReadRow;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(89[9:20])
    
    wire co_mult_10u_9u_0_0_4, mult_10u_9u_0_pp_1_10, mult_10u_9u_0_pp_1_9, 
        co_mult_10u_9u_0_0_3, mult_10u_9u_0_pp_1_8, mult_10u_9u_0_pp_1_7, 
        co_mult_10u_9u_0_0_2, mult_10u_9u_0_pp_1_6, mult_10u_9u_0_pp_1_5, 
        co_mult_10u_9u_0_0_1, mult_10u_9u_0_pp_1_4, mult_10u_9u_0_pp_1_3, 
        mult_10u_9u_0_pp_1_2, mfco_3, mult_10u_9u_0_cin_lr_6, mult_9u_9u_0_cin_lr_6, 
        mult_9u_9u_0_cin_lr_4;
    wire [7:0]SpriteRead_yInSprite_7__N_597;
    
    wire LOGIC_CLOCK_enable_13;
    wire [1:0]n2194;
    wire [7:0]xPre;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(104[9:13])
    
    wire LOGIC_CLOCK_enable_102, n3188, LOGIC_CLOCK_enable_110, mfco_2, 
        mult_10u_9u_0_cin_lr_4, mult_9u_9u_0_cin_lr_2, mfco_1, n4626, 
        mult_10u_9u_0_cin_lr_2, mult_9u_9u_0_pp_2_4, n15857, n15858;
    wire [15:0]currSprite_pos;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(191[9:23])
    
    wire n14062, n14021;
    wire [15:0]currSprite_size;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(194[9:24])
    
    wire n14022, n14061, n8_c, n14, n15728, SpriteRead_xValid_N_1167, 
        n14656;
    wire [3:0]currColor_lat;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(113[9:22])
    
    wire LOGIC_CLOCK_enable_18, n17442, n12, n15743, n14_adj_1884, 
        LOGIC_CLOCK_enable_19, LOGIC_CLOCK_enable_122;
    wire [9:0]VRAM_DATA_9__N_848;
    
    wire LOGIC_CLOCK_enable_131;
    wire [9:0]VRAM_DATA_19__N_858;
    
    wire LOGIC_CLOCK_enable_140;
    wire [9:0]VRAM_DATA_29__N_868;
    
    wire LOGIC_CLOCK_enable_157, n4485, LOGIC_CLOCK_enable_27;
    wire [15:0]n3855;
    
    wire n3960, n16082, n16083, n16086, n3935, n3936, n3937, n3938, 
        n16095, n16096, n16099, mult_9u_9u_0_cin_lr_0, mult_9u_9u_0_pp_4_16, 
        n16105, n16106, n16109, n16112, n16113, n16116, mult_9u_9u_0_pp_4_15, 
        mult_9u_9u_0_pp_4_14, mult_9u_9u_0_pp_4_13;
    wire [3:0]BUS_transferState;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(133[9:26])
    
    wire LOGIC_CLOCK_enable_48;
    wire [3:0]BUS_transferState_3__N_443;
    
    wire LOGIC_CLOCK_enable_29, n16119, n16120, n16123, n4276;
    wire [7:0]xOffset_pre;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(94[9:20])
    
    wire LOGIC_CLOCK_enable_165, n16138, n16139;
    wire [15:0]Sprite_readData2;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(174[9:25])
    
    wire LOGIC_CLOCK_enable_172, n4521, n16153, n16154, n16168, n16169, 
        n16183, n16184, n16198, n16199, n4486, MDM_done, LOGIC_CLOCK_enable_32, 
        n16213, n16214, n16228, n16229, n16249, n16250, n16253, 
        n16268, n16269, n16272, n16296, n16297, n16300, n4381, 
        n16318, n16319, n16322, n58, n62_adj_1885, n100, LOGIC_CLOCK_enable_175, 
        mult_9u_9u_0_pp_4_12, mult_9u_9u_0_pp_4_11, mult_9u_9u_0_pp_3_16, 
        mult_9u_9u_0_pp_3_15, mco_15;
    wire [14:0]Sprite_writeAddr;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(177[9:25])
    
    wire LOGIC_CLOCK_enable_196;
    wire [8:0]Sprite_writeData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(178[9:25])
    
    wire n4520, LOGIC_CLOCK_enable_38, co_mult_9u_9u_0_2_7, s_mult_9u_9u_0_1_17, 
        s_mult_9u_9u_0_2_17, mco_14, mco_13;
    wire [15:0]Sprite_readData2_15__N_492;
    wire [15:0]Sprite_readData2_15__N_476;
    
    wire mco_12, mco_11, n3955, n3956, n3957, n3958;
    wire [15:0]Sprite_readData2_15__N_524;
    wire [15:0]Sprite_readData2_15__N_508;
    
    wire mco_10, n16134, n16135, n16136, n16137, n7_c;
    wire [15:0]currSprite_conf;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(197[9:24])
    
    wire SpriteRead_yValid_N_1156;
    wire [7:0]SpriteRead_yValid_N_1158_c;
    
    wire n7_adj_1886, n46_c, n6, n16149, n16150, n16151, n16152, 
        n16164, n16165, n1193;
    wire [1:0]n898;
    
    wire n16166, n16167, n17056, n17058, mco_9, mco_8, mult_9u_9u_0_pp_2_5, 
        n16179, n16180, n16181, n16182, n16194, n16195, n16196, 
        n16197, n16209, n16210, SpriteRead_xValid_N_1166, n16772, 
        mco_7, n16211, n16212, mco_6, n16224, n16225, n16226, 
        n16227, mco_5, mco_4;
    wire [7:0]yOffset_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(97[9:16])
    
    wire n16087, n15388, n18258, mco_3_adj_1902, mco_2_adj_1903, n9918, 
        n10025, n23_adj_1904, n17283, n8626, n3198, n15444, n17433, 
        n10, n15699, n17280, n15442, n15625, n17369, n77;
    wire [7:0]n683;
    
    wire n15378, n16100, n15, mco_1_adj_1905, n16110, n15525, n17446, 
        n15375, n17460, SpriteRead_xValid, mco_adj_1906, n17406, n16773, 
        n58_adj_1908, n60, co_t_mult_9u_9u_0_3_5, n5, n17450, n16117, 
        n17268, n17485, n4416, n17459, otherData2_15__N_540, n1230, 
        n1345;
    wire [3:0]BUS_transferState_3__N_926;
    
    wire n17461, n17357, co_mult_10u_9u_0_2_5_adj_1909, s_mult_10u_9u_0_1_13_adj_1910, 
        s_mult_10u_9u_0_1_14_adj_1911, s_mult_10u_9u_0_0_13_adj_1912, s_mult_10u_9u_0_0_14_adj_1913, 
        co_mult_10u_9u_0_2_6_adj_1914, s_mult_10u_9u_0_2_13_adj_1915, s_mult_10u_9u_0_2_14_adj_1916, 
        n16124, co_mult_9u_9u_0_2_6, s_mult_9u_9u_0_1_15, s_mult_9u_9u_0_1_16, 
        s_mult_9u_9u_0_2_15, s_mult_9u_9u_0_2_16, n4310, co_mult_9u_9u_0_2_5, 
        s_mult_9u_9u_0_2_13, s_mult_9u_9u_0_2_14, n14_adj_1917, n15664, 
        n70, n2539, n4079, n4095, n16103, n4044, n4060, n16102, 
        n4188, n4076, n4092, n16093, n4153, n4172, n4057, n16092, 
        n4075, n4091, n16090, n4137, n3939, n3940, n3941, n3942, 
        n4056, n16089;
    wire [7:0]x;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(101[9:10])
    
    wire n14012, n4074, n4090, n16080, n4039, n4055, n16079, n18256, 
        n14447, n17367, n17403, n17405, n3990, n3991, n3992, n3993, 
        n15528, n17306, n16442, LOGIC_CLOCK_enable_45, co_t_mult_9u_9u_0_3_4, 
        n4073, n4089, n16077, n14153, n4038, n4054, n16076, co_mult_9u_9u_0_2_4, 
        s_mult_9u_9u_0_2_11, s_mult_9u_9u_0_2_12, s_mult_10u_9u_0_1_15_adj_1918, 
        s_mult_10u_9u_0_1_16_adj_1919, s_mult_10u_9u_0_0_15_adj_1920, co_mult_10u_9u_0_2_7_adj_1921, 
        s_mult_10u_9u_0_2_15_adj_1922, s_mult_10u_9u_0_2_16_adj_1923, s_mult_10u_9u_0_1_17_adj_1924, 
        s_mult_10u_9u_0_1_18_adj_1925, s_mult_10u_9u_0_2_17_adj_1926, s_mult_10u_9u_0_2_18_adj_1927, 
        co_mult_10u_9u_0_1_6_adj_1928, mult_10u_9u_0_pp_3_17_adj_1929, co_mult_10u_9u_0_1_5_adj_1930, 
        mult_10u_9u_0_pp_2_15_adj_1931, mult_10u_9u_0_pp_3_16_adj_1932, 
        mult_10u_9u_0_pp_3_15_adj_1933, co_mult_10u_9u_0_1_4_adj_1934, mult_10u_9u_0_pp_2_14_adj_1935, 
        mult_10u_9u_0_pp_2_13_adj_1936, mult_10u_9u_0_pp_3_14_adj_1937, 
        mult_10u_9u_0_pp_3_13_adj_1938, co_mult_10u_9u_0_1_3_adj_1939, s_mult_10u_9u_0_1_11_adj_1940, 
        s_mult_10u_9u_0_1_12_adj_1941, mult_10u_9u_0_pp_2_12_adj_1942, mult_10u_9u_0_pp_2_11_adj_1943, 
        mult_10u_9u_0_pp_3_12_adj_1944, mult_10u_9u_0_pp_3_11_adj_1945, 
        co_mult_10u_9u_0_1_2_adj_1946, s_mult_10u_9u_0_1_9_adj_1947, s_mult_10u_9u_0_1_10_adj_1948, 
        mult_10u_9u_0_pp_2_10_adj_1949, mult_10u_9u_0_pp_2_9_adj_1950, mult_10u_9u_0_pp_3_10_adj_1951, 
        mult_10u_9u_0_pp_3_9_adj_1952, co_mult_10u_9u_0_1_1_adj_1953, s_mult_10u_9u_0_1_7_adj_1954, 
        s_mult_10u_9u_0_1_8_adj_1955, mult_10u_9u_0_pp_2_8_adj_1956, mult_10u_9u_0_pp_2_7_adj_1957, 
        mult_10u_9u_0_pp_3_8_adj_1958, mult_10u_9u_0_pp_3_7_adj_1959, mult_10u_9u_0_pp_3_6_adj_1960, 
        s_mult_10u_9u_0_1_6_adj_1961, mult_10u_9u_0_pp_2_6_adj_1962, co_mult_10u_9u_0_0_7_adj_1963, 
        co_mult_10u_9u_0_0_6_adj_1964, mult_10u_9u_0_pp_1_13_adj_1965, n14060, 
        co_mult_9u_9u_0_2_3, co_mult_10u_9u_0_0_5_adj_1966, mult_10u_9u_0_pp_0_11_adj_1967, 
        s_mult_10u_9u_0_0_11_adj_1968, s_mult_10u_9u_0_0_12_adj_1969, mult_10u_9u_0_pp_1_12_adj_1970, 
        mult_10u_9u_0_pp_1_11_adj_1971, n14320, n17428, co_mult_10u_9u_0_0_4_adj_1972, 
        s_mult_10u_9u_0_0_9_adj_1973, s_mult_10u_9u_0_0_10_adj_1974, mult_10u_9u_0_pp_0_10_adj_1975, 
        mult_10u_9u_0_pp_0_9_adj_1976, mult_10u_9u_0_pp_1_10_adj_1977, mult_10u_9u_0_pp_1_9_adj_1978, 
        co_mult_9u_9u_0_1_6, n4072, n4088, n16074, ALPHA_WE, n4037, 
        n4053, n16073, n4071, n4087, n16071, n4036, n4052, n16070, 
        n17472, n4070, n4086, n16068, n4035, n4051, n16067, n4083, 
        n4084, n4085, n4069, n16065, n14152, n4093, n4094, n4048, 
        n4049, n4050, n14151, co_mult_10u_9u_0_0_3_adj_1979, s_mult_10u_9u_0_0_7_adj_1980, 
        s_mult_10u_9u_0_0_8_adj_1981, mult_10u_9u_0_pp_0_8_adj_1982, mult_10u_9u_0_pp_0_7_adj_1983, 
        mult_10u_9u_0_pp_1_8_adj_1984, mult_10u_9u_0_pp_1_7_adj_1985, n4034, 
        n16064, n14150, co_mult_10u_9u_0_0_2_adj_1986, s_mult_10u_9u_0_0_5_adj_1987, 
        s_mult_10u_9u_0_0_6_adj_1988, mult_10u_9u_0_pp_0_6_adj_1989, mult_10u_9u_0_pp_0_5_adj_1990, 
        mult_10u_9u_0_pp_1_6_adj_1991, mult_10u_9u_0_pp_1_5_adj_1992, n14149, 
        n4058, n4059;
    wire [18:0]BLUE_OUT_9__N_687;
    
    wire co_mult_10u_9u_0_0_1_adj_1993, s_mult_10u_9u_0_0_4_adj_1994, mult_10u_9u_0_pp_0_4_adj_1995, 
        mult_10u_9u_0_pp_0_3_adj_1996, mult_10u_9u_0_pp_1_4_adj_1997, mult_10u_9u_0_pp_1_3_adj_1998, 
        n4067, n4068, mult_10u_9u_0_pp_1_2_adj_1999, mult_10u_9u_0_pp_0_2_adj_2000, 
        mfco_3_adj_2001, n4077, n4078, mult_10u_9u_0_cin_lr_6_adj_2002, 
        n4032, n4033, mfco_2_adj_2003, n14148, n14147, n4080, n4081, 
        n4082, n17439;
    wire [7:0]SpriteRead_xValid_N_1168;
    
    wire n4_c, n16805, n4045, n4046, n4047, n4061, n4062, n4063, 
        n4096, n4097, n4098, n14013;
    wire [7:0]xOffset_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(96[9:16])
    
    wire n14014, n14133, n14059, LOGIC_CLOCK_enable_49, n14406, n3978, 
        n3979, n3980, n3981, n3982, n3983, n3984, n3985, n14132, 
        n3986, n3987, n3988, n3989, n14058, n6_adj_2004, n6187, 
        n14131, n3943, n3944, n3945, n3946, n17388, n14057, frameEndClock, 
        LOGIC_CLOCK_enable_50, n3947, n3948, n3949, n3950, n3951, 
        n3952, n3953, n3954, n14130, n14056;
    wire [9:0]BLUE_OUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(231[9:17])
    
    wire n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
        n3970, n3971, n3972, n3973, n3927, n3928, n3929, n3930, 
        n3931, n3932, n3933, n3934, n17451, n17468, n60_adj_2005, 
        n17429, n17443, n16062, n3974, n3975, n3976, n3977, n16061, 
        n16056, n16055, n16053, n16052, mult_10u_9u_0_cin_lr_4_adj_2006, 
        mfco_1_adj_2007, mult_10u_9u_0_cin_lr_2_adj_2008, mfco_adj_2009, 
        n16050, co_mult_9u_9u_0_2_2, mult_10u_9u_0_pp_2_4_adj_2010, mult_9u_9u_0_cin_lr_0_adj_2011, 
        mult_9u_9u_0_pp_4_16_adj_2012, mult_9u_9u_0_pp_4_15_adj_2013, mult_9u_9u_0_pp_4_14_adj_2014, 
        LOGIC_CLOCK_enable_51, Sprite_writeClk_N_1144, GR_WR_CLK_N_1081, 
        GREEN_WE, LOGIC_CLOCK_enable_53, BLUE_WE, LOGIC_CLOCK_enable_54, 
        n14129, mult_9u_9u_0_pp_4_13_adj_2015, n14055;
    wire [17:0]BLUE_OUT_9__N_706;
    
    wire mult_9u_9u_0_pp_4_12_adj_2016, mult_9u_9u_0_pp_4_11_adj_2017, mult_9u_9u_0_pp_4_10_adj_2018, 
        n14019;
    wire [7:0]y;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(102[9:10])
    
    wire n73, n17402, mult_9u_9u_0_pp_4_9_adj_2019, mult_9u_9u_0_pp_3_16_adj_2020, 
        mult_9u_9u_0_pp_3_15_adj_2021, mco_15_adj_2022, n8405, n14339, 
        n17447, n15_adj_2023, mult_9u_9u_0_pp_3_14_adj_2024, mult_9u_9u_0_pp_3_13_adj_2025, 
        mco_14_adj_2026, LOGIC_CLOCK_enable_74, mult_9u_9u_0_pp_3_12_adj_2027, 
        mult_9u_9u_0_pp_3_11_adj_2028, mco_13_adj_2029, mult_9u_9u_0_pp_3_10_adj_2030, 
        mult_9u_9u_0_pp_3_9_adj_2031, mco_12_adj_2032, mult_9u_9u_0_pp_3_8_adj_2033, 
        mult_9u_9u_0_pp_3_7_adj_2034, mult_9u_9u_0_cin_lr_6_adj_2035, mult_9u_9u_0_pp_2_14_adj_2036, 
        mult_9u_9u_0_pp_2_13_adj_2037, mco_11_adj_2038, n16049, mult_9u_9u_0_pp_2_12_adj_2039, 
        mult_9u_9u_0_pp_2_11_adj_2040, mco_10_adj_2041, co_t_mult_9u_9u_0_3_3, 
        mult_9u_9u_0_pp_2_10_adj_2042, mult_9u_9u_0_pp_2_9_adj_2043, mco_9_adj_2044, 
        n16047, n14128, n14054, n14018, n14017, mult_9u_9u_0_pp_2_8_adj_2045, 
        mult_9u_9u_0_pp_2_7_adj_2046, mco_8_adj_2047, mult_9u_9u_0_pp_2_6_adj_2048, 
        mult_9u_9u_0_pp_2_5_adj_2049, mult_9u_9u_0_cin_lr_4_adj_2050, mult_9u_9u_0_pp_1_12_adj_2051, 
        mult_9u_9u_0_pp_1_11_adj_2052, mco_7_adj_2053, mult_9u_9u_0_pp_1_10_adj_2054, 
        mult_9u_9u_0_pp_1_9_adj_2055, mco_6_adj_2056, mult_9u_9u_0_pp_1_8_adj_2057, 
        mult_9u_9u_0_pp_1_7_adj_2058, mco_5_adj_2059, mult_9u_9u_0_pp_1_6_adj_2060, 
        mult_9u_9u_0_pp_1_5_adj_2061, mco_4_adj_2062, n17349, n16046, 
        n16044, n16043, mult_9u_9u_0_pp_1_4_adj_2063, mult_9u_9u_0_pp_1_3_adj_2064, 
        mult_9u_9u_0_cin_lr_2_adj_2065, mult_9u_9u_0_pp_0_10_adj_2066, mult_9u_9u_0_pp_0_9_adj_2067, 
        mco_3_adj_2068, n14127, RED_WE, mult_9u_9u_0_pp_0_8_adj_2069, 
        mult_9u_9u_0_pp_0_7_adj_2070, mco_2_adj_2071, n17397, n14053, 
        mult_9u_9u_0_pp_0_6_adj_2072, mult_9u_9u_0_pp_0_5_adj_2073, mco_1_adj_2074, 
        n14016, n14126, n15403, n17264, n17265, n14_adj_2075, mult_9u_9u_0_pp_0_4_adj_2076, 
        mult_9u_9u_0_pp_0_3_adj_2077, mco_adj_2078;
    wire [17:0]GREEN_OUT_9__N_669;
    
    wire mult_9u_9u_0_pp_0_2_adj_2079, co_t_mult_9u_9u_0_3_5_adj_2080, s_mult_9u_9u_0_2_17_adj_2081, 
        n11, n16041, n17361, n17360, n15_adj_2082, n17263, n14052, 
        co_t_mult_9u_9u_0_3_4_adj_2083, s_mult_9u_9u_0_2_15_adj_2084, s_mult_9u_9u_0_2_16_adj_2085, 
        co_t_mult_9u_9u_0_3_3_adj_2086, s_mult_9u_9u_0_2_13_adj_2087, s_mult_9u_9u_0_2_14_adj_2088, 
        n17396, n17255, co_t_mult_9u_9u_0_3_2_adj_2089, s_mult_9u_9u_0_2_11_adj_2090, 
        s_mult_9u_9u_0_2_12_adj_2091, co_t_mult_9u_9u_0_3_1_adj_2092, s_mult_9u_9u_0_2_9_adj_2093, 
        s_mult_9u_9u_0_2_10_adj_2094, s_mult_9u_9u_0_2_8_adj_2095, co_mult_9u_9u_0_2_7_adj_2096, 
        s_mult_9u_9u_0_1_17_adj_2097;
    wire [17:0]currAddress_17__N_724;
    
    wire co_mult_9u_9u_0_2_6_adj_2098, s_mult_9u_9u_0_1_15_adj_2099, s_mult_9u_9u_0_1_16_adj_2100, 
        co_mult_9u_9u_0_2_5_adj_2101, s_mult_9u_9u_0_1_13_adj_2102, s_mult_9u_9u_0_1_14_adj_2103, 
        s_mult_9u_9u_0_0_13_adj_2104, co_mult_9u_9u_0_2_4_adj_2105, s_mult_9u_9u_0_1_11_adj_2106, 
        s_mult_9u_9u_0_1_12_adj_2107, s_mult_9u_9u_0_0_11_adj_2108, s_mult_9u_9u_0_0_12_adj_2109, 
        co_mult_9u_9u_0_2_3_adj_2110, s_mult_9u_9u_0_1_9_adj_2111, s_mult_9u_9u_0_1_10_adj_2112, 
        s_mult_9u_9u_0_0_9_adj_2113, s_mult_9u_9u_0_0_10_adj_2114, co_mult_9u_9u_0_2_2_adj_2115, 
        s_mult_9u_9u_0_1_7_adj_2116, s_mult_9u_9u_0_1_8_adj_2117, s_mult_9u_9u_0_0_7_adj_2118, 
        s_mult_9u_9u_0_0_8_adj_2119, co_mult_9u_9u_0_2_1, s_mult_9u_9u_0_1_6_adj_2120, 
        s_mult_9u_9u_0_0_5_adj_2121, s_mult_9u_9u_0_0_6_adj_2122, mult_9u_9u_0_pp_2_4_adj_2123, 
        s_mult_9u_9u_0_0_4_adj_2124, co_mult_9u_9u_0_1_6_adj_2125, co_mult_9u_9u_0_1_5_adj_2126, 
        co_mult_9u_9u_0_1_4_adj_2127, co_mult_9u_9u_0_1_3_adj_2128, n1, 
        n17271, n15701, co_mult_9u_9u_0_1_2_adj_2129, co_mult_9u_9u_0_1_1_adj_2130, 
        mult_9u_9u_0_pp_3_6_adj_2131, co_mult_9u_9u_0_0_6_adj_2132, co_mult_9u_9u_0_0_5_adj_2133, 
        co_mult_9u_9u_0_0_4_adj_2134, co_mult_9u_9u_0_0_3_adj_2135, n16040, 
        co_mult_9u_9u_0_0_2_adj_2136, co_mult_9u_9u_0_0_1_adj_2137, mult_9u_9u_0_pp_1_2_adj_2138, 
        n16038, n16037, n16035, n8625, n3201, co_mult_9u_9u_0_2_1_adj_2139, 
        mult_10u_9u_0_pp_4_8_adj_2140, n16034, n17262, n15343, n4_adj_2141, 
        mco_15_adj_2142, mco_14_adj_2143, mco_13_adj_2144, mco_12_adj_2145, 
        reset_N_1062, mco_11_adj_2146, mco_10_adj_2147, mco_9_adj_2148, 
        mco_8_adj_2149, LOGIC_CLOCK_enable_81, n14125;
    wire [13:0]n16;
    wire [15:0]Sprite_readAddr;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(180[9:24])
    
    wire n16032, n14124, n14123, mco_7_adj_2150, n17483, n17484, 
        n17318;
    wire [1:0]n2191;
    
    wire n17, n15352, mco_6_adj_2151, mco_5_adj_2152, mco_4_adj_2153, 
        n16031, co_mult_10u_9u_0_2_4_adj_2154, s_mult_10u_9u_0_2_11_adj_2155, 
        s_mult_10u_9u_0_2_12_adj_2156, co_mult_10u_9u_0_2_3_adj_2157, s_mult_10u_9u_0_2_9_adj_2158, 
        s_mult_10u_9u_0_2_10_adj_2159, co_mult_10u_9u_0_2_2_adj_2160, s_mult_10u_9u_0_2_8_adj_2161, 
        co_mult_10u_9u_0_2_1_adj_2162, mult_10u_9u_0_pp_2_5_adj_2163, co_t_mult_10u_9u_0_3_1_adj_2164, 
        mult_10u_9u_0_pp_4_9_adj_2165, mult_10u_9u_0_pp_4_10_adj_2166, co_t_mult_10u_9u_0_3_2_adj_2167, 
        mult_10u_9u_0_pp_4_11_adj_2168, mult_10u_9u_0_pp_4_12_adj_2169, 
        co_t_mult_10u_9u_0_3_3_adj_2170, mult_10u_9u_0_pp_4_13_adj_2171, 
        mult_10u_9u_0_pp_4_14_adj_2172, co_t_mult_10u_9u_0_3_4_adj_2173, 
        mult_10u_9u_0_pp_4_15_adj_2174, mult_10u_9u_0_pp_4_16_adj_2175, 
        co_t_mult_10u_9u_0_3_5_adj_2176, mult_10u_9u_0_pp_4_17_adj_2177, 
        mult_10u_9u_0_cin_lr_0_adj_2178, mco_adj_2179, mco_1_adj_2180, 
        mco_2_adj_2181, mco_3_adj_2182, mco_4_adj_2183, mco_5_adj_2184, 
        mco_6_adj_2185, mco_7_adj_2186, mco_8_adj_2187, mco_9_adj_2188, 
        mco_10_adj_2189, mco_11_adj_2190, mco_12_adj_2191, mco_13_adj_2192, 
        mco_14_adj_2193, mco_15_adj_2194, mult_9u_9u_0_pp_3_6_adj_2195, 
        mult_9u_9u_0_pp_2_4_adj_2196, mult_9u_9u_0_pp_1_2_adj_2197, mult_9u_9u_0_cin_lr_2_adj_2198, 
        mult_9u_9u_0_cin_lr_4_adj_2199, mult_9u_9u_0_cin_lr_6_adj_2200, 
        co_mult_9u_9u_0_0_1_adj_2201, mult_9u_9u_0_pp_0_2_adj_2202, co_mult_9u_9u_0_0_2_adj_2203, 
        s_mult_9u_9u_0_0_4_adj_2204, mult_9u_9u_0_pp_0_4_adj_2205, mult_9u_9u_0_pp_0_3_adj_2206, 
        mult_9u_9u_0_pp_1_4_adj_2207, mult_9u_9u_0_pp_1_3_adj_2208, co_mult_9u_9u_0_0_3_adj_2209, 
        s_mult_9u_9u_0_0_5_adj_2210, s_mult_9u_9u_0_0_6_adj_2211, mult_9u_9u_0_pp_0_6_adj_2212, 
        mult_9u_9u_0_pp_0_5_adj_2213, mult_9u_9u_0_pp_1_6_adj_2214, mult_9u_9u_0_pp_1_5_adj_2215, 
        co_mult_9u_9u_0_0_4_adj_2216, s_mult_9u_9u_0_0_7_adj_2217, s_mult_9u_9u_0_0_8_adj_2218, 
        mult_9u_9u_0_pp_0_8_adj_2219, mult_9u_9u_0_pp_0_7_adj_2220, mult_9u_9u_0_pp_1_8_adj_2221, 
        mult_9u_9u_0_pp_1_7_adj_2222, co_mult_9u_9u_0_0_5_adj_2223, s_mult_9u_9u_0_0_9_adj_2224, 
        s_mult_9u_9u_0_0_10_adj_2225, mult_9u_9u_0_pp_0_10_adj_2226, mult_9u_9u_0_pp_0_9_adj_2227, 
        mult_9u_9u_0_pp_1_10_adj_2228, mult_9u_9u_0_pp_1_9_adj_2229, co_mult_9u_9u_0_0_6_adj_2230, 
        s_mult_9u_9u_0_0_11_adj_2231, s_mult_9u_9u_0_0_12_adj_2232, mult_9u_9u_0_pp_1_12_adj_2233, 
        mult_9u_9u_0_pp_1_11_adj_2234, s_mult_9u_9u_0_0_13_adj_2235, co_mult_9u_9u_0_1_1_adj_2236, 
        s_mult_9u_9u_0_1_6_adj_2237, mult_9u_9u_0_pp_2_6_adj_2238, co_mult_9u_9u_0_1_2_adj_2239, 
        s_mult_9u_9u_0_1_7_adj_2240, s_mult_9u_9u_0_1_8_adj_2241, mult_9u_9u_0_pp_2_8_adj_2242, 
        mult_9u_9u_0_pp_2_7_adj_2243, mult_9u_9u_0_pp_3_8_adj_2244, mult_9u_9u_0_pp_3_7_adj_2245, 
        co_mult_9u_9u_0_1_3_adj_2246, s_mult_9u_9u_0_1_9_adj_2247, s_mult_9u_9u_0_1_10_adj_2248, 
        mult_9u_9u_0_pp_2_10_adj_2249, mult_9u_9u_0_pp_2_9_adj_2250, mult_9u_9u_0_pp_3_10_adj_2251, 
        mult_9u_9u_0_pp_3_9_adj_2252, co_mult_9u_9u_0_1_4_adj_2253, s_mult_9u_9u_0_1_11_adj_2254, 
        s_mult_9u_9u_0_1_12_adj_2255, mult_9u_9u_0_pp_2_12_adj_2256, mult_9u_9u_0_pp_2_11_adj_2257, 
        mult_9u_9u_0_pp_3_12_adj_2258, mult_9u_9u_0_pp_3_11_adj_2259, co_mult_9u_9u_0_1_5_adj_2260, 
        s_mult_9u_9u_0_1_13_adj_2261, s_mult_9u_9u_0_1_14_adj_2262, mult_9u_9u_0_pp_2_14_adj_2263, 
        mult_9u_9u_0_pp_2_13_adj_2264, mult_9u_9u_0_pp_3_14_adj_2265, mult_9u_9u_0_pp_3_13_adj_2266, 
        co_mult_9u_9u_0_1_6_adj_2267, s_mult_9u_9u_0_1_15_adj_2268, s_mult_9u_9u_0_1_16_adj_2269, 
        mult_9u_9u_0_pp_3_16_adj_2270, mult_9u_9u_0_pp_3_15_adj_2271, s_mult_9u_9u_0_1_17_adj_2272, 
        co_mult_9u_9u_0_2_1_adj_2273, co_mult_9u_9u_0_2_2_adj_2274, mult_9u_9u_0_pp_2_5_adj_2275, 
        co_mult_9u_9u_0_2_3_adj_2276, s_mult_9u_9u_0_2_8_adj_2277, co_mult_9u_9u_0_2_4_adj_2278, 
        s_mult_9u_9u_0_2_9_adj_2279, s_mult_9u_9u_0_2_10_adj_2280, co_mult_9u_9u_0_2_5_adj_2281, 
        s_mult_9u_9u_0_2_11_adj_2282, s_mult_9u_9u_0_2_12_adj_2283, co_mult_9u_9u_0_2_6_adj_2284, 
        s_mult_9u_9u_0_2_13_adj_2285, s_mult_9u_9u_0_2_14_adj_2286, co_mult_9u_9u_0_2_7_adj_2287, 
        s_mult_9u_9u_0_2_15_adj_2288, s_mult_9u_9u_0_2_16_adj_2289, s_mult_9u_9u_0_2_17_adj_2290, 
        co_t_mult_9u_9u_0_3_1_adj_2291, mult_9u_9u_0_pp_4_9_adj_2292, mult_9u_9u_0_pp_4_10_adj_2293, 
        co_t_mult_9u_9u_0_3_2_adj_2294, mult_9u_9u_0_pp_4_11_adj_2295, mult_9u_9u_0_pp_4_12_adj_2296, 
        co_t_mult_9u_9u_0_3_3_adj_2297, mult_9u_9u_0_pp_4_13_adj_2298, mult_9u_9u_0_pp_4_14_adj_2299, 
        co_t_mult_9u_9u_0_3_4_adj_2300, mult_9u_9u_0_pp_4_15_adj_2301, mult_9u_9u_0_pp_4_16_adj_2302, 
        co_t_mult_9u_9u_0_3_5_adj_2303, mult_9u_9u_0_cin_lr_0_adj_2304, 
        mco_adj_2305, mco_1_adj_2306, mco_2_adj_2307, mco_3_adj_2308, 
        mco_4_adj_2309, mco_5_adj_2310, mco_6_adj_2311, mco_7_adj_2312, 
        mco_8_adj_2313, mco_9_adj_2314, mco_10_adj_2315, mco_11_adj_2316, 
        mco_12_adj_2317, mco_13_adj_2318, mco_14_adj_2319, mco_15_adj_2320, 
        n16029, n16028, n16026, n5_adj_2321, n17448, n14122, n14121, 
        n16025, n14120, n14119, n15420, n17449, n15508, n16023, 
        n16022;
    wire [7:0]SpriteRead_xInSprite;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(186[9:29])
    
    wire n14051, n17404, n16020, n17257, n16019, n14050, n14049, 
        n14048, n16254, n16017, n16016, n17175, n16014, n16013, 
        n16011, n16010, n16008, n16007, n17454, n17286, n15448, 
        n16005, n16004, n5113, n16002, n14113, n14047;
    wire [9:0]GREEN_OUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(230[9:18])
    wire [3:0]BUS_transferState_3__N_930;
    
    wire n13998, n13999, n16273, n14112, n14046, n16001, n15999, 
        n15998, n15996, n14111, n15995, mult_10u_9u_0_pp_3_6_adj_2322, 
        mult_10u_9u_0_pp_2_4_adj_2323, mult_10u_9u_0_pp_1_2_adj_2324;
    wire [18:0]RED_OUT_9__N_613;
    
    wire mult_10u_9u_0_pp_0_11_adj_2325, mfco_adj_2326, mult_10u_9u_0_cin_lr_2_adj_2327, 
        mult_10u_9u_0_pp_1_13_adj_2328, mfco_1_adj_2329, mult_10u_9u_0_cin_lr_4_adj_2330, 
        mult_10u_9u_0_pp_2_15_adj_2331, mfco_2_adj_2332, mult_10u_9u_0_cin_lr_6_adj_2333, 
        mult_10u_9u_0_pp_3_17_adj_2334, mfco_3_adj_2335, co_mult_10u_9u_0_0_1_adj_2336, 
        mult_10u_9u_0_pp_0_2_adj_2337, co_mult_10u_9u_0_0_2_adj_2338, s_mult_10u_9u_0_0_4_adj_2339, 
        mult_10u_9u_0_pp_0_4_adj_2340, mult_10u_9u_0_pp_0_3_adj_2341, mult_10u_9u_0_pp_1_4_adj_2342, 
        mult_10u_9u_0_pp_1_3_adj_2343, co_mult_10u_9u_0_0_3_adj_2344, s_mult_10u_9u_0_0_5_adj_2345, 
        s_mult_10u_9u_0_0_6_adj_2346, mult_10u_9u_0_pp_0_6_adj_2347, mult_10u_9u_0_pp_0_5_adj_2348, 
        mult_10u_9u_0_pp_1_6_adj_2349, mult_10u_9u_0_pp_1_5_adj_2350, co_mult_10u_9u_0_0_4_adj_2351, 
        s_mult_10u_9u_0_0_7_adj_2352, s_mult_10u_9u_0_0_8_adj_2353, mult_10u_9u_0_pp_0_8_adj_2354, 
        mult_10u_9u_0_pp_0_7_adj_2355, mult_10u_9u_0_pp_1_8_adj_2356, mult_10u_9u_0_pp_1_7_adj_2357, 
        co_mult_10u_9u_0_0_5_adj_2358, s_mult_10u_9u_0_0_9_adj_2359, s_mult_10u_9u_0_0_10_adj_2360, 
        mult_10u_9u_0_pp_0_10_adj_2361, mult_10u_9u_0_pp_0_9_adj_2362, mult_10u_9u_0_pp_1_10_adj_2363, 
        mult_10u_9u_0_pp_1_9_adj_2364, co_mult_10u_9u_0_0_6_adj_2365, s_mult_10u_9u_0_0_11_adj_2366, 
        s_mult_10u_9u_0_0_12_adj_2367, mult_10u_9u_0_pp_1_12_adj_2368, mult_10u_9u_0_pp_1_11_adj_2369, 
        co_mult_10u_9u_0_0_7_adj_2370, s_mult_10u_9u_0_0_13_adj_2371, s_mult_10u_9u_0_0_14_adj_2372, 
        s_mult_10u_9u_0_0_15_adj_2373, co_mult_10u_9u_0_1_1_adj_2374, s_mult_10u_9u_0_1_6_adj_2375, 
        mult_10u_9u_0_pp_2_6_adj_2376, co_mult_10u_9u_0_1_2_adj_2377, s_mult_10u_9u_0_1_7_adj_2378, 
        s_mult_10u_9u_0_1_8_adj_2379, mult_10u_9u_0_pp_2_8_adj_2380, mult_10u_9u_0_pp_2_7_adj_2381, 
        mult_10u_9u_0_pp_3_8_adj_2382, mult_10u_9u_0_pp_3_7_adj_2383, co_mult_10u_9u_0_1_3_adj_2384, 
        s_mult_10u_9u_0_1_9_adj_2385, s_mult_10u_9u_0_1_10_adj_2386, mult_10u_9u_0_pp_2_10_adj_2387, 
        mult_10u_9u_0_pp_2_9_adj_2388, mult_10u_9u_0_pp_3_10_adj_2389, mult_10u_9u_0_pp_3_9_adj_2390, 
        co_mult_10u_9u_0_1_4_adj_2391, s_mult_10u_9u_0_1_11_adj_2392, s_mult_10u_9u_0_1_12_adj_2393, 
        mult_10u_9u_0_pp_2_12_adj_2394, mult_10u_9u_0_pp_2_11_adj_2395, 
        mult_10u_9u_0_pp_3_12_adj_2396, mult_10u_9u_0_pp_3_11_adj_2397, 
        co_mult_10u_9u_0_1_5_adj_2398, s_mult_10u_9u_0_1_13_adj_2399, s_mult_10u_9u_0_1_14_adj_2400, 
        mult_10u_9u_0_pp_2_14_adj_2401, mult_10u_9u_0_pp_2_13_adj_2402, 
        mult_10u_9u_0_pp_3_14_adj_2403, mult_10u_9u_0_pp_3_13_adj_2404, 
        co_mult_10u_9u_0_1_6_adj_2405, s_mult_10u_9u_0_1_15_adj_2406, s_mult_10u_9u_0_1_16_adj_2407, 
        mult_10u_9u_0_pp_3_16_adj_2408, mult_10u_9u_0_pp_3_15_adj_2409, 
        s_mult_10u_9u_0_1_17_adj_2410, s_mult_10u_9u_0_1_18_adj_2411, co_mult_10u_9u_0_2_1_adj_2412, 
        co_mult_10u_9u_0_2_2_adj_2413, mult_10u_9u_0_pp_2_5_adj_2414, co_mult_10u_9u_0_2_3_adj_2415, 
        s_mult_10u_9u_0_2_8_adj_2416, co_mult_10u_9u_0_2_4_adj_2417, s_mult_10u_9u_0_2_9_adj_2418, 
        s_mult_10u_9u_0_2_10_adj_2419, co_mult_10u_9u_0_2_5_adj_2420, s_mult_10u_9u_0_2_11_adj_2421, 
        s_mult_10u_9u_0_2_12_adj_2422, co_mult_10u_9u_0_2_6_adj_2423, s_mult_10u_9u_0_2_13_adj_2424, 
        s_mult_10u_9u_0_2_14_adj_2425, co_mult_10u_9u_0_2_7_adj_2426, s_mult_10u_9u_0_2_15_adj_2427, 
        s_mult_10u_9u_0_2_16_adj_2428, s_mult_10u_9u_0_2_17_adj_2429, s_mult_10u_9u_0_2_18_adj_2430, 
        co_t_mult_10u_9u_0_3_1_adj_2431, mult_10u_9u_0_pp_4_9_adj_2432, 
        mult_10u_9u_0_pp_4_10_adj_2433, co_t_mult_10u_9u_0_3_2_adj_2434, 
        mult_10u_9u_0_pp_4_11_adj_2435, mult_10u_9u_0_pp_4_12_adj_2436, 
        co_t_mult_10u_9u_0_3_3_adj_2437, mult_10u_9u_0_pp_4_13_adj_2438, 
        mult_10u_9u_0_pp_4_14_adj_2439, co_t_mult_10u_9u_0_3_4_adj_2440, 
        mult_10u_9u_0_pp_4_15_adj_2441, mult_10u_9u_0_pp_4_16_adj_2442, 
        co_t_mult_10u_9u_0_3_5_adj_2443, mult_10u_9u_0_pp_4_17_adj_2444, 
        mult_10u_9u_0_cin_lr_0_adj_2445, mco_adj_2446, mco_1_adj_2447, 
        mco_2_adj_2448, mco_3_adj_2449, mco_4_adj_2450, mco_5_adj_2451, 
        mco_6_adj_2452, mco_7_adj_2453, mco_8_adj_2454, mco_9_adj_2455, 
        mco_10_adj_2456, mco_11_adj_2457, mco_12_adj_2458, mco_13_adj_2459, 
        mco_14_adj_2460, mco_15_adj_2461, n14045, n3189, n3190, n3191, 
        n3192, n3193, n3194, n3195;
    wire [8:0]n949;
    
    wire LOGIC_CLOCK_enable_158, n14110, n17291, n14109, n14108, n4_adj_2464, 
        n14511, n14107, n4_adj_2465;
    wire [7:0]n30;
    
    wire n19, n15681, n21, n15457, n17284, n14106, n15689, n22_adj_2467, 
        n18, n19_adj_2468, n15693, n17180, n17179, n6135, n17480, 
        n17481, n17341, n16301, n14044, n14043, n14042, n14041, 
        n14040, n14039, n13997, n13996, n14038;
    wire [9:0]RED_OUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(229[9:16])
    
    wire n10_adj_2469, n15611, n16323, n17295, n11_adj_2470, n10_adj_2471, 
        n17297, n15725, n12_adj_2473, n15369, n14087, n14086, n14037, 
        n14085, n14036, n14084, n14002, n14035, n14083, n14034, 
        n14001, n14033, n14082, n14000, n14032, n14031, n14030, 
        n93, n14236, n14235, n17386, n15629, n14028;
    wire [7:0]n972;
    
    wire n14234, n14233, n14232, n14231, n16473, n17296, n14027, 
        n14219, n14218, n10_adj_2475;
    wire [9:0]GR_RE_DOUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(159[9:19])
    
    wire n16478, n15453, n14217, n14216, n15410, n9_adj_2477, n14215, 
        n14214, n14213, n17359, n14212, n14026, n14211, n14210, 
        n14338, n14073, n17300, n1339, n17301, n6_adj_2478, n15510, 
        n14072, n15512;
    wire [7:0]GR_WR_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(160[9:19])
    
    wire n14071, n17285, n14070, n69, n20, n14412, n13, n11_adj_2480, 
        n15714, n14069, n14068, n15635, n16632, n14023, n16771, 
        n1_adj_2481, n2, n17_adj_2482, n7044, n14067, n14066, n16058, 
        n16059, n6157, n15476, n55, n17294, n14065, n10444, n70_adj_2484, 
        n17370, n5146, n10461, n17471;
    wire [8:0]Sprite_readData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(181[9:24])
    
    MULT2 mult_10u_9u_0_mult_0_4 (.A0(VRAM_DATA_OUT[18]), .A1(VRAM_DATA_OUT[19]), 
          .A2(VRAM_DATA_OUT[19]), .A3(GND_net), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_3), .CO(mfco), .P0(mult_10u_9u_0_pp_0_9), .P1(mult_10u_9u_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_0_3 (.A0(VRAM_DATA_OUT[16]), .A1(VRAM_DATA_OUT[17]), 
          .A2(VRAM_DATA_OUT[17]), .A3(VRAM_DATA_OUT[18]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_2), .CO(mco_3), .P0(mult_10u_9u_0_pp_0_7), .P1(mult_10u_9u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    CCU2D add_617_7 (.A0(currAddress_17__N_742[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_742[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14063), .COUT(n14064), .S0(currAddress[5]), 
          .S1(currAddress[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_7.INIT0 = 16'hfaaa;
    defparam add_617_7.INIT1 = 16'hfaaa;
    defparam add_617_7.INJECT1_0 = "NO";
    defparam add_617_7.INJECT1_1 = "NO";
    MULT2 mult_10u_9u_0_mult_0_2 (.A0(VRAM_DATA_OUT[14]), .A1(VRAM_DATA_OUT[15]), 
          .A2(VRAM_DATA_OUT[15]), .A3(VRAM_DATA_OUT[16]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_1), .CO(mco_2), .P0(mult_10u_9u_0_pp_0_5), .P1(mult_10u_9u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FD1P3AX currSprite_999__i0 (.D(n37[0]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[0])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i0.GSR = "ENABLED";
    FADD2B mult_9u_9u_0_add_1_5 (.A0(mult_9u_9u_0_pp_2_13), .A1(mult_9u_9u_0_pp_2_14), 
           .B0(mult_9u_9u_0_pp_3_13), .B1(mult_9u_9u_0_pp_3_14), .CI(co_mult_9u_9u_0_1_4), 
           .COUT(co_mult_9u_9u_0_1_5), .S0(s_mult_9u_9u_0_1_13), .S1(s_mult_9u_9u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_10u_9u_0_mult_0_1 (.A0(VRAM_DATA_OUT[12]), .A1(VRAM_DATA_OUT[13]), 
          .A2(VRAM_DATA_OUT[13]), .A3(VRAM_DATA_OUT[14]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco), .CO(mco_1), .P0(mult_10u_9u_0_pp_0_3), .P1(mult_10u_9u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_0_0 (.A0(VRAM_DATA_OUT[10]), .A1(VRAM_DATA_OUT[11]), 
          .A2(VRAM_DATA_OUT[11]), .A3(VRAM_DATA_OUT[12]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mult_10u_9u_0_cin_lr_0), .CO(mco), .P0(GREEN_OUT_9__N_650[1]), 
          .P1(mult_10u_9u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B t_mult_10u_9u_0_add_3_6 (.A0(s_mult_10u_9u_0_2_17), .A1(s_mult_10u_9u_0_2_18), 
           .B0(mult_10u_9u_0_pp_4_17), .B1(GND_net), .CI(co_t_mult_10u_9u_0_3_5), 
           .S0(GREEN_OUT_9__N_650[17]), .S1(GREEN_OUT_9__N_650[18])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    PFUMX i96 (.BLUT(n59), .ALUT(n62), .C0(state[7]), .Z(n95));
    FADD2B mult_9u_9u_0_add_1_4 (.A0(mult_9u_9u_0_pp_2_11), .A1(mult_9u_9u_0_pp_2_12), 
           .B0(mult_9u_9u_0_pp_3_11), .B1(mult_9u_9u_0_pp_3_12), .CI(co_mult_9u_9u_0_1_3), 
           .COUT(co_mult_9u_9u_0_1_4), .S0(s_mult_9u_9u_0_1_11), .S1(s_mult_9u_9u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_9u_9u_0_add_1_3 (.A0(mult_9u_9u_0_pp_2_9), .A1(mult_9u_9u_0_pp_2_10), 
           .B0(mult_9u_9u_0_pp_3_9), .B1(mult_9u_9u_0_pp_3_10), .CI(co_mult_9u_9u_0_1_2), 
           .COUT(co_mult_9u_9u_0_1_3), .S0(s_mult_9u_9u_0_1_9), .S1(s_mult_9u_9u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 SRAM_WE_N_1255_I_0_269_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17382), .Z(lastAddress_31__N_1338)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_269_2_lut_3_lut_4_lut_4_lut.init = 16'hfd55;
    FADD2B mult_9u_9u_0_add_1_2 (.A0(mult_9u_9u_0_pp_2_7), .A1(mult_9u_9u_0_pp_2_8), 
           .B0(mult_9u_9u_0_pp_3_7), .B1(mult_9u_9u_0_pp_3_8), .CI(co_mult_9u_9u_0_1_1), 
           .COUT(co_mult_9u_9u_0_1_2), .S0(s_mult_9u_9u_0_1_7), .S1(s_mult_9u_9u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B t_mult_10u_9u_0_add_3_5 (.A0(s_mult_10u_9u_0_2_15), .A1(s_mult_10u_9u_0_2_16), 
           .B0(mult_10u_9u_0_pp_4_15), .B1(mult_10u_9u_0_pp_4_16), .CI(co_t_mult_10u_9u_0_3_4), 
           .COUT(co_t_mult_10u_9u_0_3_5), .S0(GREEN_OUT_9__N_650[15]), .S1(GREEN_OUT_9__N_650[16])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B Cadd_mult_9u_9u_0_1_1 (.A0(GND_net), .A1(mult_9u_9u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_9u_9u_0_1_1), 
           .S1(s_mult_9u_9u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B Cadd_mult_9u_9u_0_0_7 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_0_6), .S0(s_mult_9u_9u_0_0_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B t_mult_10u_9u_0_add_3_4 (.A0(s_mult_10u_9u_0_2_13), .A1(s_mult_10u_9u_0_2_14), 
           .B0(mult_10u_9u_0_pp_4_13), .B1(mult_10u_9u_0_pp_4_14), .CI(co_t_mult_10u_9u_0_3_3), 
           .COUT(co_t_mult_10u_9u_0_3_4), .S0(GREEN_OUT_9__N_650[13]), .S1(GREEN_OUT_9__N_650[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B t_mult_10u_9u_0_add_3_3 (.A0(s_mult_10u_9u_0_2_11), .A1(s_mult_10u_9u_0_2_12), 
           .B0(mult_10u_9u_0_pp_4_11), .B1(mult_10u_9u_0_pp_4_12), .CI(co_t_mult_10u_9u_0_3_2), 
           .COUT(co_t_mult_10u_9u_0_3_3), .S0(GREEN_OUT_9__N_650[11]), .S1(GREEN_OUT_9__N_650[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_9u_9u_0_add_0_6 (.A0(GND_net), .A1(GND_net), .B0(mult_9u_9u_0_pp_1_11), 
           .B1(mult_9u_9u_0_pp_1_12), .CI(co_mult_9u_9u_0_0_5), .COUT(co_mult_9u_9u_0_0_6), 
           .S0(s_mult_9u_9u_0_0_11), .S1(s_mult_9u_9u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B t_mult_10u_9u_0_add_3_2 (.A0(s_mult_10u_9u_0_2_9), .A1(s_mult_10u_9u_0_2_10), 
           .B0(mult_10u_9u_0_pp_4_9), .B1(mult_10u_9u_0_pp_4_10), .CI(co_t_mult_10u_9u_0_3_1), 
           .COUT(co_t_mult_10u_9u_0_3_2), .S0(GREEN_OUT_9__N_650[9]), .S1(GREEN_OUT_9__N_650[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B Cadd_t_mult_10u_9u_0_3_1 (.A0(GND_net), .A1(s_mult_10u_9u_0_2_8), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_4_8), .CI(GND_net), .COUT(co_t_mult_10u_9u_0_3_1), 
           .S1(GREEN_OUT_9__N_650[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_9u_9u_0_add_0_5 (.A0(mult_9u_9u_0_pp_0_9), .A1(mult_9u_9u_0_pp_0_10), 
           .B0(mult_9u_9u_0_pp_1_9), .B1(mult_9u_9u_0_pp_1_10), .CI(co_mult_9u_9u_0_0_4), 
           .COUT(co_mult_9u_9u_0_0_5), .S0(s_mult_9u_9u_0_0_9), .S1(s_mult_9u_9u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(s_mult_10u_9u_0_1_17), 
           .B1(s_mult_10u_9u_0_1_18), .CI(co_mult_10u_9u_0_2_7), .S0(s_mult_10u_9u_0_2_17), 
           .S1(s_mult_10u_9u_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_2_7 (.A0(s_mult_10u_9u_0_0_15), .A1(GND_net), 
           .B0(s_mult_10u_9u_0_1_15), .B1(s_mult_10u_9u_0_1_16), .CI(co_mult_10u_9u_0_2_6), 
           .COUT(co_mult_10u_9u_0_2_7), .S0(s_mult_10u_9u_0_2_15), .S1(s_mult_10u_9u_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_2_6 (.A0(s_mult_10u_9u_0_0_13), .A1(s_mult_10u_9u_0_0_14), 
           .B0(s_mult_10u_9u_0_1_13), .B1(s_mult_10u_9u_0_1_14), .CI(co_mult_10u_9u_0_2_5), 
           .COUT(co_mult_10u_9u_0_2_6), .S0(s_mult_10u_9u_0_2_13), .S1(s_mult_10u_9u_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_2_5 (.A0(s_mult_10u_9u_0_0_11), .A1(s_mult_10u_9u_0_0_12), 
           .B0(s_mult_10u_9u_0_1_11), .B1(s_mult_10u_9u_0_1_12), .CI(co_mult_10u_9u_0_2_4), 
           .COUT(co_mult_10u_9u_0_2_5), .S0(s_mult_10u_9u_0_2_11), .S1(s_mult_10u_9u_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_2_4 (.A0(s_mult_10u_9u_0_0_9), .A1(s_mult_10u_9u_0_0_10), 
           .B0(s_mult_10u_9u_0_1_9), .B1(s_mult_10u_9u_0_1_10), .CI(co_mult_10u_9u_0_2_3), 
           .COUT(co_mult_10u_9u_0_2_4), .S0(s_mult_10u_9u_0_2_9), .S1(s_mult_10u_9u_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_2_3 (.A0(s_mult_10u_9u_0_0_7), .A1(s_mult_10u_9u_0_0_8), 
           .B0(s_mult_10u_9u_0_1_7), .B1(s_mult_10u_9u_0_1_8), .CI(co_mult_10u_9u_0_2_2), 
           .COUT(co_mult_10u_9u_0_2_3), .S0(GREEN_OUT_9__N_650[7]), .S1(s_mult_10u_9u_0_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_2_2 (.A0(s_mult_10u_9u_0_0_5), .A1(s_mult_10u_9u_0_0_6), 
           .B0(mult_10u_9u_0_pp_2_5), .B1(s_mult_10u_9u_0_1_6), .CI(co_mult_10u_9u_0_2_1), 
           .COUT(co_mult_10u_9u_0_2_2), .S0(GREEN_OUT_9__N_650[5]), .S1(GREEN_OUT_9__N_650[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    LUT4 i284_2_lut (.A(LOGIC_CLOCK_enable_33), .B(lastReadRow_2_derived_5), 
         .Z(LOGIC_CLOCK_enable_113)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam i284_2_lut.init = 16'h2222;
    FADD2B Cadd_mult_10u_9u_0_2_1 (.A0(GND_net), .A1(s_mult_10u_9u_0_0_4), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_2_4), .CI(GND_net), .COUT(co_mult_10u_9u_0_2_1), 
           .S1(GREEN_OUT_9__N_650[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_1_7 (.A0(GND_net), .A1(GND_net), .B0(mult_10u_9u_0_pp_3_17), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_1_6), .S0(s_mult_10u_9u_0_1_17), 
           .S1(s_mult_10u_9u_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_9u_9u_0_add_0_4 (.A0(mult_9u_9u_0_pp_0_7), .A1(mult_9u_9u_0_pp_0_8), 
           .B0(mult_9u_9u_0_pp_1_7), .B1(mult_9u_9u_0_pp_1_8), .CI(co_mult_9u_9u_0_0_3), 
           .COUT(co_mult_9u_9u_0_0_4), .S0(s_mult_9u_9u_0_0_7), .S1(s_mult_9u_9u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FD1P3AX GR_WR_DOUT_16__i1 (.D(GR_WR_DOUT[0]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i1.GSR = "DISABLED";
    FADD2B t_mult_9u_9u_0_add_3_2 (.A0(s_mult_9u_9u_0_2_9), .A1(s_mult_9u_9u_0_2_10), 
           .B0(mult_9u_9u_0_pp_4_9), .B1(mult_9u_9u_0_pp_4_10), .CI(co_t_mult_9u_9u_0_3_1), 
           .COUT(co_t_mult_9u_9u_0_3_2), .S0(RED_OUT_9__N_632[9]), .S1(RED_OUT_9__N_632[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_9u_9u_0_add_0_3 (.A0(mult_9u_9u_0_pp_0_5), .A1(mult_9u_9u_0_pp_0_6), 
           .B0(mult_9u_9u_0_pp_1_5), .B1(mult_9u_9u_0_pp_1_6), .CI(co_mult_9u_9u_0_0_2), 
           .COUT(co_mult_9u_9u_0_0_3), .S0(s_mult_9u_9u_0_0_5), .S1(s_mult_9u_9u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_add_1_6 (.A0(mult_10u_9u_0_pp_2_15), .A1(GND_net), 
           .B0(mult_10u_9u_0_pp_3_15), .B1(mult_10u_9u_0_pp_3_16), .CI(co_mult_10u_9u_0_1_5), 
           .COUT(co_mult_10u_9u_0_1_6), .S0(s_mult_10u_9u_0_1_15), .S1(s_mult_10u_9u_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_1_5 (.A0(mult_10u_9u_0_pp_2_13), .A1(mult_10u_9u_0_pp_2_14), 
           .B0(mult_10u_9u_0_pp_3_13), .B1(mult_10u_9u_0_pp_3_14), .CI(co_mult_10u_9u_0_1_4), 
           .COUT(co_mult_10u_9u_0_1_5), .S0(s_mult_10u_9u_0_1_13), .S1(s_mult_10u_9u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    PFUMX mux_634_i8 (.BLUT(otherData[7]), .ALUT(n2872[7]), .C0(n1985), 
          .Z(\BUS_DATA_INTERNAL[7] ));
    FD1S3AX yOffset_i0 (.D(yOffset_pre[0]), .CK(offsetLatchClockOrd), .Q(yOffset[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i0.GSR = "DISABLED";
    DPR16X4C Sprite_sizes4 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4380), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4040), .DO1(n4041), .DO2(n4042), .DO3(n4043));
    defparam Sprite_sizes4.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d02 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4311), 
            .DO0(n4305), .DO1(n4306), .DO2(n4307), .DO3(n4308));
    defparam Sprite_positions_d02.initval = "0x0000000000000000";
    AND2 AND2_t8 (.A(RED_READ[0]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(167[10:63])
    FADD2B Cadd_t_mult_9u_9u_0_3_1 (.A0(GND_net), .A1(s_mult_9u_9u_0_2_8), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_4_8), .CI(GND_net), .COUT(co_t_mult_9u_9u_0_3_1), 
           .S1(RED_OUT_9__N_632[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_add_1_4 (.A0(mult_10u_9u_0_pp_2_11), .A1(mult_10u_9u_0_pp_2_12), 
           .B0(mult_10u_9u_0_pp_3_11), .B1(mult_10u_9u_0_pp_3_12), .CI(co_mult_10u_9u_0_1_3), 
           .COUT(co_mult_10u_9u_0_1_4), .S0(s_mult_10u_9u_0_1_11), .S1(s_mult_10u_9u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FD1S3AX state_i0 (.D(state_7__N_336[0]), .CK(LOGIC_CLOCK), .Q(\state[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i0.GSR = "ENABLED";
    AND2 AND2_t9 (.A(VRAM_DATA_OUT[10]), .B(RED_OUT_9__N_768[8]), .Z(mult_10u_9u_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(178[10:64])
    AND2 AND2_t8_adj_278 (.A(GREEN_READ[0]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_8_adj_1880)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(167[10:63])
    PFUMX mux_634_i7 (.BLUT(otherData[6]), .ALUT(n2872[6]), .C0(n1985), 
          .Z(\BUS_DATA_INTERNAL[6] ));
    AND2 AND2_t9_adj_279 (.A(VRAM_DATA_OUT[20]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_8_adj_1881)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(178[10:64])
    AND2 AND2_t8_adj_280 (.A(BLUE_READ[0]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_8_adj_1882)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(167[10:63])
    FADD2B mult_10u_9u_0_add_1_3 (.A0(mult_10u_9u_0_pp_2_9), .A1(mult_10u_9u_0_pp_2_10), 
           .B0(mult_10u_9u_0_pp_3_9), .B1(mult_10u_9u_0_pp_3_10), .CI(co_mult_10u_9u_0_1_2), 
           .COUT(co_mult_10u_9u_0_1_3), .S0(s_mult_10u_9u_0_1_9), .S1(s_mult_10u_9u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FD1P3DX latchForce_729 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_4), 
            .CK(LOGIC_CLOCK), .CD(n17276), .Q(latchForce)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam latchForce_729.GSR = "DISABLED";
    FADD2B mult_10u_9u_0_add_1_2 (.A0(mult_10u_9u_0_pp_2_7), .A1(mult_10u_9u_0_pp_2_8), 
           .B0(mult_10u_9u_0_pp_3_7), .B1(mult_10u_9u_0_pp_3_8), .CI(co_mult_10u_9u_0_1_1), 
           .COUT(co_mult_10u_9u_0_1_2), .S0(s_mult_10u_9u_0_1_7), .S1(s_mult_10u_9u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_9u_9u_0_add_0_2 (.A0(mult_9u_9u_0_pp_0_3), .A1(mult_9u_9u_0_pp_0_4), 
           .B0(mult_9u_9u_0_pp_1_3), .B1(mult_9u_9u_0_pp_1_4), .CI(co_mult_9u_9u_0_0_1), 
           .COUT(co_mult_9u_9u_0_0_2), .S0(RED_OUT_9__N_632[3]), .S1(s_mult_9u_9u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B Cadd_mult_10u_9u_0_1_1 (.A0(GND_net), .A1(mult_10u_9u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_10u_9u_0_1_1), 
           .S1(s_mult_10u_9u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B Cadd_mult_10u_9u_0_0_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_0_7), .S0(s_mult_10u_9u_0_0_15)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_0_7 (.A0(GND_net), .A1(GND_net), .B0(mult_10u_9u_0_pp_1_13), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_0_6), .COUT(co_mult_10u_9u_0_0_7), 
           .S0(s_mult_10u_9u_0_0_13), .S1(s_mult_10u_9u_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FD1P3AX currValue_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i0.GSR = "DISABLED";
    LUT4 GR_WR_DOUT_16_15__I_0_i1_3_lut (.A(GR_WR_DOUT_16[0]), .B(otherData2[0]), 
         .C(n17314), .Z(otherData[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i1_3_lut.init = 16'hcaca;
    FADD2B mult_10u_9u_0_add_0_6 (.A0(mult_10u_9u_0_pp_0_11), .A1(GND_net), 
           .B0(mult_10u_9u_0_pp_1_11), .B1(mult_10u_9u_0_pp_1_12), .CI(co_mult_10u_9u_0_0_5), 
           .COUT(co_mult_10u_9u_0_0_6), .S0(s_mult_10u_9u_0_0_11), .S1(s_mult_10u_9u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B Cadd_mult_9u_9u_0_0_1 (.A0(GND_net), .A1(mult_9u_9u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_9u_9u_0_0_1), 
           .S1(RED_OUT_9__N_632[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FD1P3IX currColor_998__i3 (.D(n3[3]), .SP(LOGIC_CLOCK_enable_33), .CD(n7210), 
            .CK(LOGIC_CLOCK), .Q(currColor[3]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_998__i3.GSR = "ENABLED";
    FD1P3IX currColor_998__i2 (.D(n3[2]), .SP(LOGIC_CLOCK_enable_33), .CD(n7210), 
            .CK(LOGIC_CLOCK), .Q(currColor[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_998__i2.GSR = "ENABLED";
    FD1P3IX currColor_998__i1 (.D(n3[1]), .SP(LOGIC_CLOCK_enable_33), .CD(n7210), 
            .CK(LOGIC_CLOCK), .Q(currColor[1]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_998__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n17334), .B(n17321), .C(n17273), .D(n17312), 
         .Z(n4415)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(577[24:69])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    PFUMX mux_634_i6 (.BLUT(otherData[5]), .ALUT(n2872[5]), .C0(n1985), 
          .Z(\BUS_DATA_INTERNAL[5] ));
    FD1S1A currReadRow_4__I_0_798_i1 (.D(\SpriteRead_yInSprite_7__N_597[0] ), 
           .CK(lastReadRow_2_derived_5), .Q(lastReadRow[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(294[2] 453[14])
    defparam currReadRow_4__I_0_798_i1.GSR = "DISABLED";
    FADD2B mult_10u_9u_0_add_0_5 (.A0(mult_10u_9u_0_pp_0_9), .A1(mult_10u_9u_0_pp_0_10), 
           .B0(mult_10u_9u_0_pp_1_9), .B1(mult_10u_9u_0_pp_1_10), .CI(co_mult_10u_9u_0_0_4), 
           .COUT(co_mult_10u_9u_0_0_5), .S0(s_mult_10u_9u_0_0_9), .S1(s_mult_10u_9u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_0_4 (.A0(mult_10u_9u_0_pp_0_7), .A1(mult_10u_9u_0_pp_0_8), 
           .B0(mult_10u_9u_0_pp_1_7), .B1(mult_10u_9u_0_pp_1_8), .CI(co_mult_10u_9u_0_0_3), 
           .COUT(co_mult_10u_9u_0_0_4), .S0(s_mult_10u_9u_0_0_7), .S1(s_mult_10u_9u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_0_3 (.A0(mult_10u_9u_0_pp_0_5), .A1(mult_10u_9u_0_pp_0_6), 
           .B0(mult_10u_9u_0_pp_1_5), .B1(mult_10u_9u_0_pp_1_6), .CI(co_mult_10u_9u_0_0_2), 
           .COUT(co_mult_10u_9u_0_0_3), .S0(s_mult_10u_9u_0_0_5), .S1(s_mult_10u_9u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_add_0_2 (.A0(mult_10u_9u_0_pp_0_3), .A1(mult_10u_9u_0_pp_0_4), 
           .B0(mult_10u_9u_0_pp_1_3), .B1(mult_10u_9u_0_pp_1_4), .CI(co_mult_10u_9u_0_0_1), 
           .COUT(co_mult_10u_9u_0_0_2), .S0(GREEN_OUT_9__N_650[3]), .S1(s_mult_10u_9u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B Cadd_mult_10u_9u_0_0_1 (.A0(GND_net), .A1(mult_10u_9u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_10u_9u_0_0_1), 
           .S1(GREEN_OUT_9__N_650[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_Cadd_6_5 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(mult_10u_9u_0_pp_3_17)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_9u_9u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_9u_9u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FD1P3AX currRowOffset__i1 (.D(n2194[0]), .SP(LOGIC_CLOCK_enable_13), 
            .CK(LOGIC_CLOCK), .Q(SpriteRead_yInSprite_7__N_597[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currRowOffset__i1.GSR = "ENABLED";
    FD1P3AX xPre__i0 (.D(n3188), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i0.GSR = "ENABLED";
    FD1P3AX VRAM_ADDR__i1 (.D(SpriteRead_yInSprite_7__N_597[5]), .SP(LOGIC_CLOCK_enable_110), 
            .CK(LOGIC_CLOCK), .Q(\VRAM_ADDR[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i1.GSR = "DISABLED";
    FADD2B mult_10u_9u_0_Cadd_4_5 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(mult_10u_9u_0_pp_2_15)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_10u_9u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FADD2B mult_9u_9u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_Cadd_2_5 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(mult_10u_9u_0_pp_1_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    PFUMX mux_634_i5 (.BLUT(otherData[4]), .ALUT(n2872[4]), .C0(n1985), 
          .Z(\BUS_DATA_INTERNAL[4] ));
    SPR16X4C Sprite_pointers_d315 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4626), 
            .DO0(n4608), .DO1(n4609), .DO2(n4610), .DO3(n4611));
    defparam Sprite_pointers_d315.initval = "0x0000000000000000";
    SPR16X4C Sprite_pointers_d314 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4626), 
            .DO0(n4612), .DO1(n4613), .DO2(n4614), .DO3(n4615));
    defparam Sprite_pointers_d314.initval = "0x0000000000000000";
    SPR16X4C Sprite_pointers_d313 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4626), 
            .DO0(n4616), .DO1(n4617), .DO2(n4618), .DO3(n4619));
    defparam Sprite_pointers_d313.initval = "0x0000000000000000";
    FADD2B mult_10u_9u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    SPR16X4C Sprite_pointers_d312 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4591), 
            .DO0(n4573), .DO1(n4574), .DO2(n4575), .DO3(n4576));
    defparam Sprite_pointers_d312.initval = "0x0000000000000000";
    FADD2B mult_10u_9u_0_Cadd_0_5 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(mult_10u_9u_0_pp_0_11)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    LUT4 SRAM_WE_N_1255_I_0_254_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17381), .Z(lastAddress_31__N_1323)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_254_2_lut_3_lut_4_lut_4_lut.init = 16'hfd55;
    SPR16X4C Sprite_pointers_d311 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4591), 
            .DO0(n4577), .DO1(n4578), .DO2(n4579), .DO3(n4580));
    defparam Sprite_pointers_d311.initval = "0x0000000000000000";
    AND2 AND2_t12 (.A(RED_READ[0]), .B(ALPHA_READ[0]), .Z(RED_OUT_9__N_632[0])) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(159[10:64])
    SPR16X4C Sprite_pointers_d310 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4591), 
            .DO0(n4581), .DO1(n4582), .DO2(n4583), .DO3(n4584));
    defparam Sprite_pointers_d310.initval = "0x0000000000000000";
    SPR16X4C Sprite_pointers_d39 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4625), 
            .DO0(n4592), .DO1(n4593), .DO2(n4594), .DO3(n4595));
    defparam Sprite_pointers_d39.initval = "0x0000000000000000";
    AND2 AND2_t11 (.A(RED_READ[0]), .B(ALPHA_READ[2]), .Z(mult_9u_9u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(161[10:64])
    SPR16X4C Sprite_pointers_d38 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4625), 
            .DO0(n4596), .DO1(n4597), .DO2(n4598), .DO3(n4599));
    defparam Sprite_pointers_d38.initval = "0x0000000000000000";
    AND2 AND2_t10 (.A(RED_READ[0]), .B(ALPHA_READ[4]), .Z(mult_9u_9u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(163[10:64])
    SPR16X4C Sprite_pointers_d37 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4625), 
            .DO0(n4600), .DO1(n4601), .DO2(n4602), .DO3(n4603));
    defparam Sprite_pointers_d37.initval = "0x0000000000000000";
    PFUMX mux_634_i4 (.BLUT(otherData[3]), .ALUT(n2877), .C0(n1985), .Z(\BUS_DATA_INTERNAL[3] ));
    SPR16X4C Sprite_pointers_d36 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4590), 
            .DO0(n4557), .DO1(n4558), .DO2(n4559), .DO3(n4560));
    defparam Sprite_pointers_d36.initval = "0x0000000000000000";
    PFUMX i12197 (.BLUT(n15857), .ALUT(n15858), .C0(currSprite[5]), .Z(currSprite_pos[6]));
    SPR16X4C Sprite_pointers_d35 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4590), 
            .DO0(n4561), .DO1(n4562), .DO2(n4563), .DO3(n4564));
    defparam Sprite_pointers_d35.initval = "0x0000000000000000";
    AND2 AND2_t9_adj_281 (.A(RED_READ[0]), .B(ALPHA_READ[6]), .Z(mult_9u_9u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(165[10:63])
    LUT4 SRAM_WE_N_1255_I_0_297_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17373), .D(n18270), .Z(lastAddress_31__N_1413)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_297_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    PFUMX mux_634_i3 (.BLUT(otherData[2]), .ALUT(n2878), .C0(n1985), .Z(\BUS_DATA_INTERNAL[2] ));
    CCU2D add_617_5 (.A0(currColor[3]), .B0(currAddress_17__N_742[3]), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_742[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14062), .COUT(n14063), .S0(currAddress[3]), 
          .S1(currAddress[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_5.INIT0 = 16'h5666;
    defparam add_617_5.INIT1 = 16'hfaaa;
    defparam add_617_5.INJECT1_0 = "NO";
    defparam add_617_5.INJECT1_1 = "NO";
    PFUMX mux_634_i2 (.BLUT(otherData[1]), .ALUT(n2879), .C0(n1985), .Z(\BUS_DATA_INTERNAL[1] ));
    CCU2D add_19_4 (.A0(currSprite_pos[10]), .B0(currSprite_size[10]), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[11]), .B1(currSprite_size[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14021), .COUT(n14022), .S0(SpriteRead_yValid_N_1158[2]), 
          .S1(SpriteRead_yValid_N_1158[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[132:154])
    defparam add_19_4.INIT0 = 16'h5666;
    defparam add_19_4.INIT1 = 16'h5666;
    defparam add_19_4.INJECT1_0 = "NO";
    defparam add_19_4.INJECT1_1 = "NO";
    PFUMX mux_634_i1 (.BLUT(otherData[0]), .ALUT(n2880), .C0(n1985), .Z(\BUS_DATA_INTERNAL[0] ));
    CCU2D add_617_3 (.A0(currColor[1]), .B0(currAddress_17__N_742[1]), .C0(GND_net), 
          .D0(GND_net), .A1(currColor[2]), .B1(currAddress_17__N_742[2]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14061), .COUT(n14062), .S0(currAddress[1]), 
          .S1(currAddress[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_3.INIT0 = 16'h5666;
    defparam add_617_3.INIT1 = 16'h5666;
    defparam add_617_3.INJECT1_0 = "NO";
    defparam add_617_3.INJECT1_1 = "NO";
    SPR16X4C Sprite_pointers_d30 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4625), 
            .DO0(n4604), .DO1(n4605), .DO2(n4606), .DO3(n4607));
    defparam Sprite_pointers_d30.initval = "0x0000000000000000";
    PFUMX xPre_7__I_0_i16 (.BLUT(n8_c), .ALUT(n14), .C0(n15728), .Z(SpriteRead_xValid_N_1167)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;
    FD1S3AX VRAM_WC_696 (.D(n14656), .CK(LOGIC_CLOCK), .Q(VRAM_WC)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_WC_696.GSR = "ENABLED";
    FD1P3AX currColor_lat_i0_i0 (.D(currColor[0]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currColor_lat_i0_i0.GSR = "DISABLED";
    FD1P3AX Sprite_readClk_702 (.D(n17442), .SP(LOGIC_CLOCK_enable_18), 
            .CK(LOGIC_CLOCK), .Q(Sprite_readClk)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam Sprite_readClk_702.GSR = "ENABLED";
    PFUMX SpriteRead_yInSprite_7__N_597_7__I_0_i14 (.BLUT(n8), .ALUT(n12), 
          .C0(n15743), .Z(n14_adj_1884)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;
    FD1P3AX SpriteLut_readClk_703 (.D(\state[0] ), .SP(LOGIC_CLOCK_enable_19), 
            .CK(LOGIC_CLOCK), .Q(SpriteLut_readClk)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam SpriteLut_readClk_703.GSR = "ENABLED";
    FD1P3AX data_0___i1 (.D(VRAM_DATA_9__N_848[0]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i1.GSR = "DISABLED";
    FD1P3AX data_1___i1 (.D(VRAM_DATA_19__N_858[0]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i1.GSR = "DISABLED";
    FD1P3AX data_2___i1 (.D(VRAM_DATA_29__N_868[0]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[20])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i1.GSR = "DISABLED";
    AND2 AND2_t13 (.A(VRAM_DATA_OUT[10]), .B(RED_OUT_9__N_768[0]), .Z(GREEN_OUT_9__N_650[0])) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(170[10:65])
    FD1P3AX BUS_ADDR_INTERNAL__i1 (.D(currAddress[0]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i1.GSR = "DISABLED";
    SPR16X4C Sprite_sizes_d14 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4380), .DO0(n4355), 
            .DO1(n4356), .DO2(n4357), .DO3(n4358));
    defparam Sprite_sizes_d14.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d24 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4485), .DO0(n4460), 
            .DO1(n4461), .DO2(n4462), .DO3(n4463));
    defparam Sprite_options_d24.initval = "0x0000000000000000";
    SPR16X4C Sprite_pointers_d34 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4590), 
            .DO0(n4565), .DO1(n4566), .DO2(n4567), .DO3(n4568));
    defparam Sprite_pointers_d34.initval = "0x0000000000000000";
    AND2 AND2_t12_adj_282 (.A(VRAM_DATA_OUT[10]), .B(RED_OUT_9__N_768[2]), 
         .Z(mult_10u_9u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(172[10:65])
    AND2 AND2_t11_adj_283 (.A(VRAM_DATA_OUT[10]), .B(RED_OUT_9__N_768[4]), 
         .Z(mult_10u_9u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(174[10:65])
    AND2 AND2_t10_adj_284 (.A(VRAM_DATA_OUT[10]), .B(RED_OUT_9__N_768[6]), 
         .Z(mult_10u_9u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(176[10:65])
    PDPW8KC Sprite_pointers0 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .DI4(BUS_data[4]), .DI5(BUS_data[5]), .DI6(BUS_data[6]), 
            .DI7(BUS_data[7]), .DI8(BUS_data[8]), .DI9(BUS_data[9]), .DI10(BUS_data[10]), 
            .DI11(BUS_data[11]), .DI12(BUS_data[12]), .DI13(BUS_data[13]), 
            .DI14(BUS_data[14]), .DI15(BUS_data[15]), .DI16(GND_net), 
            .DI17(GND_net), .ADW0(n17339), .ADW1(n17333), .ADW2(n17332), 
            .ADW3(n17331), .ADW4(n17321), .ADW5(n17334), .ADW6(GND_net), 
            .ADW7(GND_net), .ADW8(GND_net), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(Sprite_pointers_N_1123), .CLKW(LOGIC_CLOCK), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(currSprite[0]), .ADR5(currSprite[1]), 
            .ADR6(currSprite[2]), .ADR7(currSprite[3]), .ADR8(currSprite[4]), 
            .ADR9(currSprite[5]), .ADR10(GND_net), .ADR11(GND_net), .ADR12(GND_net), 
            .CER(LOGIC_CLOCK_enable_27), .OCER(VCC_net), .CLKR(LOGIC_CLOCK), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(n3855[9]), .DO1(n3855[10]), .DO2(n3855[11]), .DO3(n3855[12]), 
            .DO4(n3855[13]), .DO9(n3855[0]), .DO10(n3855[1]), .DO11(n3855[2]), 
            .DO12(n3855[3]), .DO13(n3855[4]), .DO14(n3855[5]), .DO15(n3855[6]), 
            .DO16(n3855[7]), .DO17(n3855[8]));
    defparam Sprite_pointers0.DATA_WIDTH_W = 18;
    defparam Sprite_pointers0.DATA_WIDTH_R = 18;
    defparam Sprite_pointers0.REGMODE = "NOREG";
    defparam Sprite_pointers0.CSDECODE_W = "0b000";
    defparam Sprite_pointers0.CSDECODE_R = "0b000";
    defparam Sprite_pointers0.GSR = "DISABLED";
    defparam Sprite_pointers0.RESETMODE = "SYNC";
    defparam Sprite_pointers0.ASYNC_RESET_RELEASE = "SYNC";
    defparam Sprite_pointers0.INIT_DATA = "STATIC";
    defparam Sprite_pointers0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam Sprite_pointers0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    SPR16X4C Sprite_positions_d04 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n3960), 
            .DO0(n4250), .DO1(n4251), .DO2(n4252), .DO3(n4253));
    defparam Sprite_positions_d04.initval = "0x0000000000000000";
    L6MUX21 i12424 (.D0(n16082), .D1(n16083), .SD(n17342), .Z(n16086));
    DPR16X4C Sprite_positions4 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n3960), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3935), .DO1(n3936), .DO2(n3937), .DO3(n3938));
    defparam Sprite_positions4.initval = "0x0000000000000000";
    L6MUX21 i12437 (.D0(n16095), .D1(n16096), .SD(n17342), .Z(n16099));
    FADD2B mult_9u_9u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    AND2 AND2_t0 (.A(RED_READ[8]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(183[10:64])
    L6MUX21 i12447 (.D0(n16105), .D1(n16106), .SD(n17342), .Z(n16109));
    L6MUX21 i12454 (.D0(n16112), .D1(n16113), .SD(n17342), .Z(n16116));
    AND2 AND2_t1 (.A(RED_READ[7]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_15)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(181[10:64])
    AND2 AND2_t2 (.A(RED_READ[6]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(179[10:64])
    AND2 AND2_t3 (.A(RED_READ[5]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_13)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(177[10:64])
    FD1P3DX BUS_transferState_i1 (.D(BUS_transferState_3__N_443[1]), .SP(LOGIC_CLOCK_enable_48), 
            .CK(LOGIC_CLOCK), .CD(n17276), .Q(BUS_transferState[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam BUS_transferState_i1.GSR = "DISABLED";
    FD1P3AX currRowOffset__i2 (.D(n2194[1]), .SP(LOGIC_CLOCK_enable_29), 
            .CK(LOGIC_CLOCK), .Q(SpriteRead_yInSprite_7__N_597[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currRowOffset__i2.GSR = "ENABLED";
    L6MUX21 i12461 (.D0(n16119), .D1(n16120), .SD(n17342), .Z(n16123));
    LUT4 i1_2_lut_3_lut_4_lut_adj_285 (.A(n17321), .B(n17334), .C(n17273), 
         .D(n17310), .Z(n4276)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(573[21:66])
    defparam i1_2_lut_3_lut_4_lut_adj_285.init = 16'h0020;
    SPR16X4C Sprite_pointers_d33 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4590), 
            .DO0(n4569), .DO1(n4570), .DO2(n4571), .DO3(n4572));
    defparam Sprite_pointers_d33.initval = "0x0000000000000000";
    FD1P3AX xOffset_pre_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i0.GSR = "DISABLED";
    L6MUX21 i12478 (.D0(n16138), .D1(n16139), .SD(n17342), .Z(Sprite_readData2[9]));
    FD1P3AX yOffset_pre_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i0.GSR = "DISABLED";
    SPR16X4C Sprite_pointers_d31 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4591), 
            .DO0(n4585), .DO1(n4586), .DO2(n4587), .DO3(n4588));
    defparam Sprite_pointers_d31.initval = "0x0000000000000000";
    SPR16X4C Sprite_pointers_d32 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4626), 
            .DO0(n4620), .DO1(n4621), .DO2(n4622), .DO3(n4623));
    defparam Sprite_pointers_d32.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d215 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4521), 
            .DO0(n4503), .DO1(n4504), .DO2(n4505), .DO3(n4506));
    defparam Sprite_options_d215.initval = "0x0000000000000000";
    L6MUX21 i12493 (.D0(n16153), .D1(n16154), .SD(n17342), .Z(\Sprite_readData2[10] ));
    SPR16X4C Sprite_options_d214 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4521), 
            .DO0(n4507), .DO1(n4508), .DO2(n4509), .DO3(n4510));
    defparam Sprite_options_d214.initval = "0x0000000000000000";
    LUT4 SRAM_WE_N_1255_I_0_268_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17371), .D(n18270), .Z(lastAddress_31__N_1337)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_268_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    L6MUX21 i12508 (.D0(n16168), .D1(n16169), .SD(n17342), .Z(\Sprite_readData2[11] ));
    L6MUX21 i12523 (.D0(n16183), .D1(n16184), .SD(n17342), .Z(\Sprite_readData2[12] ));
    L6MUX21 i12538 (.D0(n16198), .D1(n16199), .SD(n17342), .Z(\Sprite_readData2[13] ));
    SPR16X4C Sprite_options_d213 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4521), 
            .DO0(n4511), .DO1(n4512), .DO2(n4513), .DO3(n4514));
    defparam Sprite_options_d213.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d212 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4486), 
            .DO0(n4468), .DO1(n4469), .DO2(n4470), .DO3(n4471));
    defparam Sprite_options_d212.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d211 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4486), 
            .DO0(n4472), .DO1(n4473), .DO2(n4474), .DO3(n4475));
    defparam Sprite_options_d211.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d210 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4486), 
            .DO0(n4476), .DO1(n4477), .DO2(n4478), .DO3(n4479));
    defparam Sprite_options_d210.initval = "0x0000000000000000";
    FD1P3DX transferDone_727 (.D(n18280), .SP(LOGIC_CLOCK_enable_32), .CK(LOGIC_CLOCK), 
            .CD(n17276), .Q(MDM_done)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam transferDone_727.GSR = "DISABLED";
    L6MUX21 i12553 (.D0(n16213), .D1(n16214), .SD(n17342), .Z(\Sprite_readData2[14] ));
    FD1P3IX currColor_998__i0 (.D(n3[0]), .SP(LOGIC_CLOCK_enable_33), .CD(n7210), 
            .CK(LOGIC_CLOCK), .Q(currColor[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_998__i0.GSR = "ENABLED";
    L6MUX21 i12568 (.D0(n16228), .D1(n16229), .SD(n17342), .Z(\Sprite_readData2[15] ));
    L6MUX21 i12591 (.D0(n16249), .D1(n16250), .SD(n17342), .Z(n16253));
    L6MUX21 i12610 (.D0(n16268), .D1(n16269), .SD(n17342), .Z(n16272));
    L6MUX21 i12638 (.D0(n16296), .D1(n16297), .SD(n17342), .Z(n16300));
    LUT4 i1_2_lut_3_lut_4_lut_adj_286 (.A(n17321), .B(n17334), .C(n17273), 
         .D(n17312), .Z(n4381)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(573[21:66])
    defparam i1_2_lut_3_lut_4_lut_adj_286.init = 16'h0020;
    L6MUX21 i12660 (.D0(n16318), .D1(n16319), .SD(n17342), .Z(n16322));
    PFUMX i101 (.BLUT(n58), .ALUT(n62_adj_1885), .C0(state[7]), .Z(n100));
    FD1P3AX latchMode_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(latchMode[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam latchMode_i0_i0.GSR = "DISABLED";
    AND2 AND2_t4 (.A(RED_READ[4]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(175[10:64])
    AND2 AND2_t5 (.A(RED_READ[3]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_11)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(173[10:64])
    AND2 AND2_t6 (.A(RED_READ[2]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(171[10:64])
    AND2 AND2_t7 (.A(RED_READ[1]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_9)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(169[10:63])
    MULT2 mult_9u_9u_0_mult_6_4 (.A0(RED_READ[8]), .A1(GND_net), .A2(GND_net), 
          .A3(GND_net), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), 
          .B3(ALPHA_READ[6]), .CI(mco_15), .P0(mult_9u_9u_0_pp_3_15), 
          .P1(mult_9u_9u_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FD1P3AX Sprite_writeAddr__i1 (.D(n17343), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i1.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i0.GSR = "DISABLED";
    SPR16X4C Sprite_options_d29 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4520), .DO0(n4487), 
            .DO1(n4488), .DO2(n4489), .DO3(n4490));
    defparam Sprite_options_d29.initval = "0x0000000000000000";
    FD1S3AX xOffset_i0 (.D(xOffset_pre[0]), .CK(offsetLatchClockOrd), .Q(xOffset[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i0.GSR = "DISABLED";
    FD1P3AY VRAM_WE_705 (.D(\state[1] ), .SP(LOGIC_CLOCK_enable_38), .CK(LOGIC_CLOCK), 
            .Q(VRAM_WE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_WE_705.GSR = "ENABLED";
    FADD2B mult_9u_9u_0_add_2_8 (.A0(GND_net), .A1(GND_net), .B0(s_mult_9u_9u_0_1_17), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_2_7), .S0(s_mult_9u_9u_0_2_17)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_6_3 (.A0(RED_READ[6]), .A1(RED_READ[7]), .A2(RED_READ[7]), 
          .A3(RED_READ[8]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), 
          .B3(ALPHA_READ[6]), .CI(mco_14), .CO(mco_15), .P0(mult_9u_9u_0_pp_3_13), 
          .P1(mult_9u_9u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_6_2 (.A0(RED_READ[4]), .A1(RED_READ[5]), .A2(RED_READ[5]), 
          .A3(RED_READ[6]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), 
          .B3(ALPHA_READ[6]), .CI(mco_13), .CO(mco_14), .P0(mult_9u_9u_0_pp_3_11), 
          .P1(mult_9u_9u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    L6MUX21 i12421 (.D0(Sprite_readData2_15__N_492[5]), .D1(Sprite_readData2_15__N_476[5]), 
            .SD(n17343), .Z(n16083));
    MULT2 mult_9u_9u_0_mult_6_1 (.A0(RED_READ[2]), .A1(RED_READ[3]), .A2(RED_READ[3]), 
          .A3(RED_READ[4]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), 
          .B3(ALPHA_READ[6]), .CI(mco_12), .CO(mco_13), .P0(mult_9u_9u_0_pp_3_9), 
          .P1(mult_9u_9u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_6_0 (.A0(RED_READ[0]), .A1(RED_READ[1]), .A2(RED_READ[1]), 
          .A3(RED_READ[2]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), 
          .B3(ALPHA_READ[6]), .CI(mult_9u_9u_0_cin_lr_6), .CO(mco_12), 
          .P0(mult_9u_9u_0_pp_3_7), .P1(mult_9u_9u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_4_4 (.A0(RED_READ[8]), .A1(GND_net), .A2(GND_net), 
          .A3(GND_net), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), 
          .B3(ALPHA_READ[4]), .CI(mco_11), .P0(mult_9u_9u_0_pp_2_13), 
          .P1(mult_9u_9u_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    SPR16X4C Sprite_options_d28 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4520), .DO0(n4491), 
            .DO1(n4492), .DO2(n4493), .DO3(n4494));
    defparam Sprite_options_d28.initval = "0x0000000000000000";
    L6MUX21 i12434 (.D0(Sprite_readData2_15__N_492[1]), .D1(Sprite_readData2_15__N_476[1]), 
            .SD(n17343), .Z(n16096));
    SPR16X4C Sprite_options_d27 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4520), .DO0(n4495), 
            .DO1(n4496), .DO2(n4497), .DO3(n4498));
    defparam Sprite_options_d27.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d26 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4485), .DO0(n4452), 
            .DO1(n4453), .DO2(n4454), .DO3(n4455));
    defparam Sprite_options_d26.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions1 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), 
            .WAD2(n17332), .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4276), 
            .RAD0(currSprite[0]), .RAD1(currSprite[1]), .RAD2(currSprite[2]), 
            .RAD3(currSprite[3]), .DO0(n3955), .DO1(n3956), .DO2(n3957), 
            .DO3(n3958));
    defparam Sprite_positions1.initval = "0x0000000000000000";
    L6MUX21 i12444 (.D0(Sprite_readData2_15__N_492[6]), .D1(Sprite_readData2_15__N_476[6]), 
            .SD(n17343), .Z(n16106));
    L6MUX21 i12450 (.D0(Sprite_readData2_15__N_524[7]), .D1(Sprite_readData2_15__N_508[7]), 
            .SD(n17343), .Z(n16112));
    L6MUX21 i12451 (.D0(Sprite_readData2_15__N_492[7]), .D1(Sprite_readData2_15__N_476[7]), 
            .SD(n17343), .Z(n16113));
    L6MUX21 i12457 (.D0(Sprite_readData2_15__N_524[8]), .D1(Sprite_readData2_15__N_508[8]), 
            .SD(n17343), .Z(n16119));
    MULT2 mult_9u_9u_0_mult_4_3 (.A0(RED_READ[6]), .A1(RED_READ[7]), .A2(RED_READ[7]), 
          .A3(RED_READ[8]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), 
          .B3(ALPHA_READ[4]), .CI(mco_10), .CO(mco_11), .P0(mult_9u_9u_0_pp_2_11), 
          .P1(mult_9u_9u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    L6MUX21 i12458 (.D0(Sprite_readData2_15__N_492[8]), .D1(Sprite_readData2_15__N_476[8]), 
            .SD(n17343), .Z(n16120));
    L6MUX21 i12656 (.D0(Sprite_readData2_15__N_524[4]), .D1(Sprite_readData2_15__N_508[4]), 
            .SD(n17343), .Z(n16318));
    L6MUX21 i12634 (.D0(Sprite_readData2_15__N_524[3]), .D1(Sprite_readData2_15__N_508[3]), 
            .SD(n17343), .Z(n16296));
    L6MUX21 i12476 (.D0(n16134), .D1(n16135), .SD(n17343), .Z(n16138));
    L6MUX21 i12477 (.D0(n16136), .D1(n16137), .SD(n17343), .Z(n16139));
    LUT4 i2_4_lut (.A(lastReadRow[3]), .B(lastReadRow[0]), .C(n17366), 
         .D(MATRIX_CURRROW[0]), .Z(n7_c)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)))+!A (B (C+(D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[11:36])
    defparam i2_4_lut.init = 16'hde7b;
    LUT4 i2_3_lut_4_lut (.A(currSprite_conf[0]), .B(SpriteRead_yValid_N_1156), 
         .C(n14_adj_1884), .D(SpriteRead_yValid_N_1158_c[7]), .Z(n7_adj_1886)) /* synthesis lut_function=(!((B (C+(D)))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h222a;
    LUT4 PIC_addr_31__I_0_i4_2_lut_rep_363_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[3] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[3]_adj_2 ), 
         .Z(n17371)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;
    defparam PIC_addr_31__I_0_i4_2_lut_rep_363_3_lut_4_lut_4_lut.init = 16'h2c20;
    LUT4 i1_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[3] ), .B(\BUS_currGrantID[0] ), 
         .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[3]_adj_2 ), .Z(n46_c)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B)) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd3df;
    LUT4 i1_4_lut (.A(lastReadRow[1]), .B(lastReadRow[4]), .C(n17453), 
         .D(n17326), .Z(n6)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[11:36])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 PIC_addr_31__I_0_i15_3_lut_rep_375_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[14] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[14]_adj_3 ), 
         .Z(n17383)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i15_3_lut_rep_375_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i3_3_lut_rep_374_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[2] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[2]_adj_4 ), 
         .Z(n17382)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i3_3_lut_rep_374_4_lut_4_lut.init = 16'h3808;
    L6MUX21 i12491 (.D0(n16149), .D1(n16150), .SD(n17343), .Z(n16153));
    L6MUX21 i12492 (.D0(n16151), .D1(n16152), .SD(n17343), .Z(n16154));
    LUT4 i1_3_lut_rep_373_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[17] ), .B(\BUS_currGrantID[0] ), 
         .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[17]_adj_5 ), .Z(n17381)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam i1_3_lut_rep_373_4_lut_4_lut.init = 16'h3808;
    LUT4 i2_2_lut_rep_264_3_lut_3_lut (.A(n17276), .B(n1985), .C(n18260), 
         .Z(n17272)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(458[95:155])
    defparam i2_2_lut_rep_264_3_lut_3_lut.init = 16'hefef;
    LUT4 PIC_addr_31__I_0_i6_3_lut_rep_372_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[5] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[5]_adj_6 ), 
         .Z(n17380)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i6_3_lut_rep_372_4_lut_4_lut.init = 16'h3808;
    L6MUX21 i12506 (.D0(n16164), .D1(n16165), .SD(n17343), .Z(n16168));
    SPR16X4C Sprite_options_d25 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4485), .DO0(n4456), 
            .DO1(n4457), .DO2(n4458), .DO3(n4459));
    defparam Sprite_options_d25.initval = "0x0000000000000000";
    LUT4 i6570_2_lut (.A(SpriteRead_yInSprite_7__N_597[5]), .B(n1193), .Z(n898[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(383[6] 396[13])
    defparam i6570_2_lut.init = 16'h4444;
    FD1S3AX state_i7 (.D(state_7__N_336[7]), .CK(LOGIC_CLOCK), .Q(state[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i7.GSR = "ENABLED";
    L6MUX21 i12507 (.D0(n16166), .D1(n16167), .SD(n17343), .Z(n16169));
    L6MUX21 i12606 (.D0(Sprite_readData2_15__N_524[2]), .D1(Sprite_readData2_15__N_508[2]), 
            .SD(n17343), .Z(n16268));
    LUT4 PIC_addr_31__I_0_i14_3_lut_rep_371_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[13] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[13]_adj_7 ), 
         .Z(n17379)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i14_3_lut_rep_371_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i9_3_lut_rep_370_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[8] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[8]_adj_8 ), 
         .Z(n17378)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i9_3_lut_rep_370_4_lut_4_lut.init = 16'h3808;
    LUT4 LED_c_bdd_2_lut_13351_3_lut (.A(n17056), .B(\state[0] ), .C(\state[1] ), 
         .Z(n17058)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam LED_c_bdd_2_lut_13351_3_lut.init = 16'h8080;
    L6MUX21 i12587 (.D0(Sprite_readData2_15__N_524[0]), .D1(Sprite_readData2_15__N_508[0]), 
            .SD(n17343), .Z(n16249));
    MULT2 mult_9u_9u_0_mult_4_2 (.A0(RED_READ[4]), .A1(RED_READ[5]), .A2(RED_READ[5]), 
          .A3(RED_READ[6]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), 
          .B3(ALPHA_READ[4]), .CI(mco_9), .CO(mco_10), .P0(mult_9u_9u_0_pp_2_9), 
          .P1(mult_9u_9u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_4_1 (.A0(RED_READ[2]), .A1(RED_READ[3]), .A2(RED_READ[3]), 
          .A3(RED_READ[4]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), 
          .B3(ALPHA_READ[4]), .CI(mco_8), .CO(mco_9), .P0(mult_9u_9u_0_pp_2_7), 
          .P1(mult_9u_9u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 PIC_addr_31__I_0_i10_3_lut_rep_368_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[9] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[9]_adj_9 ), 
         .Z(n17376)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i10_3_lut_rep_368_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i5_3_lut_rep_367_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[4] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[4]_adj_10 ), 
         .Z(n17375)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i5_3_lut_rep_367_4_lut_4_lut.init = 16'h3808;
    MULT2 mult_9u_9u_0_mult_4_0 (.A0(RED_READ[0]), .A1(RED_READ[1]), .A2(RED_READ[1]), 
          .A3(RED_READ[2]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), 
          .B3(ALPHA_READ[4]), .CI(mult_9u_9u_0_cin_lr_4), .CO(mco_8), 
          .P0(mult_9u_9u_0_pp_2_5), .P1(mult_9u_9u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 i1_3_lut_4_lut_4_lut_adj_287 (.A(n17275), .B(\state[1]_adj_11 ), 
         .C(n17434), .D(n17457), .Z(n15469)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_287.init = 16'h3020;
    L6MUX21 i12521 (.D0(n16179), .D1(n16180), .SD(n17343), .Z(n16183));
    LUT4 PIC_addr_31__I_0_i7_3_lut_rep_366_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[6] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[6]_adj_12 ), 
         .Z(n17374)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i7_3_lut_rep_366_4_lut_4_lut.init = 16'h3808;
    L6MUX21 i12522 (.D0(n16181), .D1(n16182), .SD(n17343), .Z(n16184));
    L6MUX21 i12536 (.D0(n16194), .D1(n16195), .SD(n17343), .Z(n16198));
    LUT4 PIC_addr_31__I_0_i8_3_lut_rep_365_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[7] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[7]_adj_13 ), 
         .Z(n17373)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i8_3_lut_rep_365_4_lut_4_lut.init = 16'h3808;
    L6MUX21 i12537 (.D0(n16196), .D1(n16197), .SD(n17343), .Z(n16199));
    L6MUX21 i12551 (.D0(n16209), .D1(n16210), .SD(n17343), .Z(n16213));
    LUT4 n14447_bdd_3_lut_4_lut (.A(\state[0] ), .B(state[4]), .C(SpriteRead_xValid_N_1166), 
         .D(SpriteRead_xValid_N_1167), .Z(n16772)) /* synthesis lut_function=(!(A+(B (C (D))))) */ ;
    defparam n14447_bdd_3_lut_4_lut.init = 16'h1555;
    LUT4 PIC_addr_31__I_0_i13_3_lut_rep_369_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[12] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[12]_adj_14 ), 
         .Z(n17377)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i13_3_lut_rep_369_4_lut_4_lut.init = 16'h3808;
    MULT2 mult_9u_9u_0_mult_2_4 (.A0(RED_READ[8]), .A1(GND_net), .A2(GND_net), 
          .A3(GND_net), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), 
          .B3(ALPHA_READ[2]), .CI(mco_7), .P0(mult_9u_9u_0_pp_1_11), .P1(mult_9u_9u_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    L6MUX21 i12552 (.D0(n16211), .D1(n16212), .SD(n17343), .Z(n16214));
    MULT2 mult_9u_9u_0_mult_2_3 (.A0(RED_READ[6]), .A1(RED_READ[7]), .A2(RED_READ[7]), 
          .A3(RED_READ[8]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), 
          .B3(ALPHA_READ[2]), .CI(mco_6), .CO(mco_7), .P0(mult_9u_9u_0_pp_1_9), 
          .P1(mult_9u_9u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    L6MUX21 i12566 (.D0(n16224), .D1(n16225), .SD(n17343), .Z(n16228));
    L6MUX21 i12567 (.D0(n16226), .D1(n16227), .SD(n17343), .Z(n16229));
    MULT2 mult_9u_9u_0_mult_2_2 (.A0(RED_READ[4]), .A1(RED_READ[5]), .A2(RED_READ[5]), 
          .A3(RED_READ[6]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), 
          .B3(ALPHA_READ[2]), .CI(mco_5), .CO(mco_6), .P0(mult_9u_9u_0_pp_1_7), 
          .P1(mult_9u_9u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    L6MUX21 i12588 (.D0(Sprite_readData2_15__N_492[0]), .D1(Sprite_readData2_15__N_476[0]), 
            .SD(n17343), .Z(n16250));
    LUT4 i6888_2_lut_rep_325_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[3]_adj_2 ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[3] ), 
         .Z(n17333)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam i6888_2_lut_rep_325_3_lut_4_lut_4_lut.init = 16'h3b0b;
    L6MUX21 i12607 (.D0(Sprite_readData2_15__N_492[2]), .D1(Sprite_readData2_15__N_476[2]), 
            .SD(n17343), .Z(n16269));
    FD1S1A currReadRow_4__I_0_798_i2 (.D(n17453), .CK(lastReadRow_2_derived_5), 
           .Q(lastReadRow[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(294[2] 453[14])
    defparam currReadRow_4__I_0_798_i2.GSR = "DISABLED";
    FD1S1A currReadRow_4__I_0_798_i3 (.D(n17407), .CK(lastReadRow_2_derived_5), 
           .Q(lastReadRow[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(294[2] 453[14])
    defparam currReadRow_4__I_0_798_i3.GSR = "DISABLED";
    FD1S1A currReadRow_4__I_0_798_i4 (.D(n17366), .CK(lastReadRow_2_derived_5), 
           .Q(lastReadRow[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(294[2] 453[14])
    defparam currReadRow_4__I_0_798_i4.GSR = "DISABLED";
    FD1S1A currReadRow_4__I_0_798_i5 (.D(n17326), .CK(lastReadRow_2_derived_5), 
           .Q(lastReadRow[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(294[2] 453[14])
    defparam currReadRow_4__I_0_798_i5.GSR = "DISABLED";
    L6MUX21 i12443 (.D0(Sprite_readData2_15__N_524[6]), .D1(Sprite_readData2_15__N_508[6]), 
            .SD(n17343), .Z(n16105));
    L6MUX21 i12433 (.D0(Sprite_readData2_15__N_524[1]), .D1(Sprite_readData2_15__N_508[1]), 
            .SD(n17343), .Z(n16095));
    LUT4 PIC_addr_31__I_0_i17_3_lut_rep_354_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[16] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[16]_adj_15 ), 
         .Z(n17362)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i17_3_lut_rep_354_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i16_3_lut_rep_347_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[15] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[15]_adj_16 ), 
         .Z(n17355)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i16_3_lut_rep_347_4_lut_4_lut.init = 16'h3808;
    L6MUX21 i12420 (.D0(Sprite_readData2_15__N_524[5]), .D1(Sprite_readData2_15__N_508[5]), 
            .SD(n17343), .Z(n16082));
    MULT2 mult_9u_9u_0_mult_2_1 (.A0(RED_READ[2]), .A1(RED_READ[3]), .A2(RED_READ[3]), 
          .A3(RED_READ[4]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), 
          .B3(ALPHA_READ[2]), .CI(mco_4), .CO(mco_5), .P0(mult_9u_9u_0_pp_1_5), 
          .P1(mult_9u_9u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FD1S3AX state_i6 (.D(state_7__N_336[6]), .CK(LOGIC_CLOCK), .Q(state[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i6.GSR = "ENABLED";
    FD1S3AX state_i5 (.D(state_7__N_336[5]), .CK(LOGIC_CLOCK), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i5.GSR = "ENABLED";
    FD1S3AX state_i4 (.D(state_7__N_336[4]), .CK(LOGIC_CLOCK), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i4.GSR = "ENABLED";
    FD1S3AX state_i3 (.D(state_7__N_336[3]), .CK(LOGIC_CLOCK), .Q(\state[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i3.GSR = "ENABLED";
    FD1S3AX state_i2 (.D(state_7__N_336[2]), .CK(LOGIC_CLOCK), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(state_7__N_336[1]), .CK(LOGIC_CLOCK), .Q(\state[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam state_i1.GSR = "ENABLED";
    FD1S3AX yOffset_i7 (.D(yOffset_pre[7]), .CK(offsetLatchClockOrd), .Q(yOffset_c[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i7.GSR = "DISABLED";
    FD1S3AX yOffset_i6 (.D(yOffset_pre[6]), .CK(offsetLatchClockOrd), .Q(yOffset_c[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i6.GSR = "DISABLED";
    FD1S3AX yOffset_i5 (.D(yOffset_pre[5]), .CK(offsetLatchClockOrd), .Q(yOffset_c[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i5.GSR = "DISABLED";
    FD1S3AX yOffset_i4 (.D(yOffset_pre[4]), .CK(offsetLatchClockOrd), .Q(yOffset_c[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i4.GSR = "DISABLED";
    FD1S3AX yOffset_i3 (.D(yOffset_pre[3]), .CK(offsetLatchClockOrd), .Q(\yOffset[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i3.GSR = "DISABLED";
    FD1S3AX yOffset_i2 (.D(yOffset_pre[2]), .CK(offsetLatchClockOrd), .Q(\yOffset[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i2.GSR = "DISABLED";
    FD1S3AX yOffset_i1 (.D(yOffset_pre[1]), .CK(offsetLatchClockOrd), .Q(\yOffset[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam yOffset_i1.GSR = "DISABLED";
    L6MUX21 i12635 (.D0(Sprite_readData2_15__N_492[3]), .D1(Sprite_readData2_15__N_476[3]), 
            .SD(n17343), .Z(n16297));
    L6MUX21 i12657 (.D0(Sprite_readData2_15__N_492[4]), .D1(Sprite_readData2_15__N_476[4]), 
            .SD(n17343), .Z(n16319));
    PFUMX i12425 (.BLUT(n16084), .ALUT(n16085), .C0(n17342), .Z(n16087));
    SPR16X4C Sprite_options_d20 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4520), 
            .DO0(n4499), .DO1(n4500), .DO2(n4501), .DO3(n4502));
    defparam Sprite_options_d20.initval = "0x0000000000000000";
    LUT4 i1_4_lut_adj_288 (.A(state[7]), .B(state[6]), .C(n15388), .D(n18258), 
         .Z(state_7__N_336[6])) /* synthesis lut_function=(A (B+!(C))+!A !((D)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_adj_288.init = 16'h8ace;
    MULT2 mult_9u_9u_0_mult_2_0 (.A0(RED_READ[0]), .A1(RED_READ[1]), .A2(RED_READ[1]), 
          .A3(RED_READ[2]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), 
          .B3(ALPHA_READ[2]), .CI(mult_9u_9u_0_cin_lr_2), .CO(mco_4), 
          .P0(mult_9u_9u_0_pp_1_3), .P1(mult_9u_9u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_0_4 (.A0(RED_READ[8]), .A1(GND_net), .A2(GND_net), 
          .A3(GND_net), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), 
          .B3(ALPHA_READ[0]), .CI(mco_3_adj_1902), .P0(mult_9u_9u_0_pp_0_9), 
          .P1(mult_9u_9u_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_0_3 (.A0(RED_READ[6]), .A1(RED_READ[7]), .A2(RED_READ[7]), 
          .A3(RED_READ[8]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), 
          .B3(ALPHA_READ[0]), .CI(mco_2_adj_1903), .CO(mco_3_adj_1902), 
          .P0(mult_9u_9u_0_pp_0_7), .P1(mult_9u_9u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 i1_4_lut_adj_289 (.A(state[5]), .B(\state[3] ), .C(n9918), .D(n10025), 
         .Z(n15388)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_289.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_290 (.A(SpriteRead_yValid_N_1156), .B(n14_adj_1884), 
         .C(SpriteRead_yValid_N_1158_c[7]), .D(currSprite_conf[0]), .Z(n23_adj_1904)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[32:254])
    defparam i1_2_lut_3_lut_4_lut_adj_290.init = 16'ha800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_291 (.A(SpriteRead_yValid_N_1156), .B(n14_adj_1884), 
         .C(SpriteRead_yValid_N_1158_c[7]), .D(currSprite_conf[0]), .Z(n1193)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[32:254])
    defparam i1_2_lut_3_lut_4_lut_adj_291.init = 16'h5700;
    LUT4 SpriteRead_yValid_I_0_2_lut_rep_275_3_lut (.A(SpriteRead_yValid_N_1156), 
         .B(n14_adj_1884), .C(SpriteRead_yValid_N_1158_c[7]), .Z(n17283)) /* synthesis lut_function=(A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[32:254])
    defparam SpriteRead_yValid_I_0_2_lut_rep_275_3_lut.init = 16'ha8a8;
    LUT4 i5283_3_lut_3_lut_4_lut (.A(SpriteRead_xValid_N_1166), .B(SpriteRead_xValid_N_1167), 
         .C(state[4]), .D(n8626), .Z(n3198)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i5283_3_lut_3_lut_4_lut.init = 16'h7f70;
    LUT4 i1_4_lut_adj_292 (.A(n15444), .B(state[5]), .C(n17433), .D(n10), 
         .Z(state_7__N_336[5])) /* synthesis lut_function=(A+(B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_adj_292.init = 16'heeae;
    LUT4 i3_4_lut (.A(n15699), .B(n17280), .C(state[2]), .D(n15442), 
         .Z(n15444)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i3_4_lut.init = 16'h0100;
    LUT4 i70_3_lut_rep_272_4_lut (.A(n23_adj_1904), .B(SpriteRead_xValid_N_1166), 
         .C(SpriteRead_xValid_N_1167), .D(state[4]), .Z(n17280)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i70_3_lut_rep_272_4_lut.init = 16'hc0aa;
    LUT4 i5061_4_lut_4_lut (.A(\state[3] ), .B(state[2]), .C(state[4]), 
         .D(\state[1] ), .Z(n15625)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(87[9:14])
    defparam i5061_4_lut_4_lut.init = 16'h1808;
    LUT4 i2_4_lut_adj_293 (.A(\state[0] ), .B(n17369), .C(n77), .D(n683[4]), 
         .Z(n15378)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i2_4_lut_adj_293.init = 16'hfcfe;
    PFUMX i12438 (.BLUT(n16097), .ALUT(n16098), .C0(n17342), .Z(n16100));
    LUT4 i1_3_lut (.A(state[2]), .B(\state[0] ), .C(n15), .Z(n77)) /* synthesis lut_function=(A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_3_lut.init = 16'ha8a8;
    LUT4 i6575_2_lut (.A(state[4]), .B(n17275), .Z(n683[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(320[5] 347[12])
    defparam i6575_2_lut.init = 16'h8888;
    MULT2 mult_9u_9u_0_mult_0_2 (.A0(RED_READ[4]), .A1(RED_READ[5]), .A2(RED_READ[5]), 
          .A3(RED_READ[6]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), 
          .B3(ALPHA_READ[0]), .CI(mco_1_adj_1905), .CO(mco_2_adj_1903), 
          .P0(mult_9u_9u_0_pp_0_5), .P1(mult_9u_9u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    PFUMX i12448 (.BLUT(n16107), .ALUT(n16108), .C0(n17342), .Z(n16110));
    LUT4 i12981_4_lut (.A(\state[3] ), .B(state[2]), .C(n15525), .D(n17058), 
         .Z(state_7__N_336[3])) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i12981_4_lut.init = 16'h23af;
    LUT4 i3_4_lut_adj_294 (.A(n17446), .B(n15375), .C(state[2]), .D(n17460), 
         .Z(n15525)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i3_4_lut_adj_294.init = 16'hfffd;
    LUT4 i1_4_lut_adj_295 (.A(state[7]), .B(state[4]), .C(n33), .D(SpriteRead_xValid), 
         .Z(n15375)) /* synthesis lut_function=(A (B (D))+!A (B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_adj_295.init = 16'hcd45;
    MULT2 mult_9u_9u_0_mult_0_1 (.A0(RED_READ[2]), .A1(RED_READ[3]), .A2(RED_READ[3]), 
          .A3(RED_READ[4]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), 
          .B3(ALPHA_READ[0]), .CI(mco_adj_1906), .CO(mco_1_adj_1905), 
          .P0(mult_9u_9u_0_pp_0_3), .P1(mult_9u_9u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_0_0 (.A0(RED_READ[0]), .A1(RED_READ[1]), .A2(RED_READ[1]), 
          .A3(RED_READ[2]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), 
          .B3(ALPHA_READ[0]), .CI(mult_9u_9u_0_cin_lr_0), .CO(mco_adj_1906), 
          .P0(RED_OUT_9__N_632[1]), .P1(mult_9u_9u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 PIC_addr_31__I_0_i1_3_lut_rep_377_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[0] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[0]_adj_17 ), 
         .Z(n17385)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam PIC_addr_31__I_0_i1_3_lut_rep_377_4_lut_4_lut.init = 16'h3808;
    LUT4 i12996_4_lut (.A(state[2]), .B(n100), .C(n17406), .D(n16773), 
         .Z(state_7__N_336[2])) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i12996_4_lut.init = 16'h3222;
    LUT4 i13036_3_lut (.A(n58_adj_1908), .B(\state[0] ), .C(n60), .Z(state_7__N_336[1])) /* synthesis lut_function=(!(A+(B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i13036_3_lut.init = 16'h1515;
    FADD2B t_mult_9u_9u_0_add_3_6 (.A0(s_mult_9u_9u_0_2_17), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(co_t_mult_9u_9u_0_3_5), .S0(RED_OUT_9__N_632[17])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 i1_4_lut_adj_296 (.A(\state[1] ), .B(n5), .C(n17446), .D(n17450), 
         .Z(n58_adj_1908)) /* synthesis lut_function=(!(A+!(B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_adj_296.init = 16'h5545;
    PFUMX i12455 (.BLUT(n16114), .ALUT(n16115), .C0(n17342), .Z(n16117));
    SPR16X4C Sprite_options_d23 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4485), 
            .DO0(n4464), .DO1(n4465), .DO2(n4466), .DO3(n4467));
    defparam Sprite_options_d23.initval = "0x0000000000000000";
    SPR16X4C Sprite_options_d21 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4486), 
            .DO0(n4480), .DO1(n4481), .DO2(n4482), .DO3(n4483));
    defparam Sprite_options_d21.initval = "0x0000000000000000";
    LUT4 i83_4_lut (.A(n17268), .B(n17446), .C(state[7]), .D(n15625), 
         .Z(n60)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i83_4_lut.init = 16'hca0a;
    SPR16X4C Sprite_options_d22 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4521), 
            .DO0(n4515), .DO1(n4516), .DO2(n4517), .DO3(n4518));
    defparam Sprite_options_d22.initval = "0x0000000000000000";
    LUT4 i1_4_lut_adj_297 (.A(state[7]), .B(n17485), .C(state[4]), .D(n9891), 
         .Z(n5)) /* synthesis lut_function=(A (B)+!A (B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_adj_297.init = 16'hdcdd;
    SPR16X4C Sprite_sizes_d115 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4416), .DO0(n4398), 
            .DO1(n4399), .DO2(n4400), .DO3(n4401));
    defparam Sprite_sizes_d115.initval = "0x0000000000000000";
    LUT4 i301_2_lut_3_lut_4_lut (.A(BUS_transferState[2]), .B(n17459), .C(otherData2_15__N_540), 
         .D(BUS_DONE_OUT_N_1051), .Z(n1230)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(565[8:32])
    defparam i301_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 BUS_transferState_3__I_0_779_i2_3_lut_4_lut (.A(BUS_transferState[2]), 
         .B(n17459), .C(n1345), .D(BUS_transferState_3__N_926[1]), .Z(BUS_transferState_3__N_443[1])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(565[8:32])
    defparam BUS_transferState_3__I_0_779_i2_3_lut_4_lut.init = 16'hefe0;
    SPR16X4C Sprite_sizes_d114 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4416), .DO0(n4402), 
            .DO1(n4403), .DO2(n4404), .DO3(n4405));
    defparam Sprite_sizes_d114.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d113 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4416), .DO0(n4406), 
            .DO1(n4407), .DO2(n4408), .DO3(n4409));
    defparam Sprite_sizes_d113.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d112 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4381), .DO0(n4363), 
            .DO1(n4364), .DO2(n4365), .DO3(n4366));
    defparam Sprite_sizes_d112.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d111 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4381), .DO0(n4367), 
            .DO1(n4368), .DO2(n4369), .DO3(n4370));
    defparam Sprite_sizes_d111.initval = "0x0000000000000000";
    LUT4 i3_3_lut_rep_349_4_lut (.A(state[5]), .B(n17461), .C(state[4]), 
         .D(n15442), .Z(n17357)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i3_3_lut_rep_349_4_lut.init = 16'h1000;
    FADD2B mult_10u_9u_0_add_2_6_adj_298 (.A0(s_mult_10u_9u_0_0_13_adj_1912), 
           .A1(s_mult_10u_9u_0_0_14_adj_1913), .B0(s_mult_10u_9u_0_1_13_adj_1910), 
           .B1(s_mult_10u_9u_0_1_14_adj_1911), .CI(co_mult_10u_9u_0_2_5_adj_1909), 
           .COUT(co_mult_10u_9u_0_2_6_adj_1914), .S0(s_mult_10u_9u_0_2_13_adj_1915), 
           .S1(s_mult_10u_9u_0_2_14_adj_1916)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    SPR16X4C Sprite_sizes_d110 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4381), .DO0(n4371), 
            .DO1(n4372), .DO2(n4373), .DO3(n4374));
    defparam Sprite_sizes_d110.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d19 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4415), .DO0(n4382), 
            .DO1(n4383), .DO2(n4384), .DO3(n4385));
    defparam Sprite_sizes_d19.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d18 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4415), .DO0(n4386), 
            .DO1(n4387), .DO2(n4388), .DO3(n4389));
    defparam Sprite_sizes_d18.initval = "0x0000000000000000";
    PFUMX i12462 (.BLUT(n16121), .ALUT(n16122), .C0(n17342), .Z(n16124));
    SPR16X4C Sprite_sizes_d17 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4415), .DO0(n4390), 
            .DO1(n4391), .DO2(n4392), .DO3(n4393));
    defparam Sprite_sizes_d17.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d16 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4380), .DO0(n4347), 
            .DO1(n4348), .DO2(n4349), .DO3(n4350));
    defparam Sprite_sizes_d16.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d15 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4380), .DO0(n4351), 
            .DO1(n4352), .DO2(n4353), .DO3(n4354));
    defparam Sprite_sizes_d15.initval = "0x0000000000000000";
    PFUMX i12472 (.BLUT(n16126), .ALUT(n16127), .C0(n17334), .Z(n16134));
    FADD2B mult_9u_9u_0_add_2_7 (.A0(GND_net), .A1(GND_net), .B0(s_mult_9u_9u_0_1_15), 
           .B1(s_mult_9u_9u_0_1_16), .CI(co_mult_9u_9u_0_2_6), .COUT(co_mult_9u_9u_0_2_7), 
           .S0(s_mult_9u_9u_0_2_15), .S1(s_mult_9u_9u_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    PFUMX i12473 (.BLUT(n16128), .ALUT(n16129), .C0(n17334), .Z(n16135));
    PFUMX i12474 (.BLUT(n16130), .ALUT(n16131), .C0(n17334), .Z(n16136));
    SPR16X4C Sprite_sizes_d10 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4415), .DO0(n4394), 
            .DO1(n4395), .DO2(n4396), .DO3(n4397));
    defparam Sprite_sizes_d10.initval = "0x0000000000000000";
    PFUMX i12475 (.BLUT(n16132), .ALUT(n16133), .C0(n17334), .Z(n16137));
    SPR16X4C Sprite_sizes_d13 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4380), .DO0(n4359), 
            .DO1(n4360), .DO2(n4361), .DO3(n4362));
    defparam Sprite_sizes_d13.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes_d11 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4381), .DO0(n4375), 
            .DO1(n4376), .DO2(n4377), .DO3(n4378));
    defparam Sprite_sizes_d11.initval = "0x0000000000000000";
    LUT4 i1_2_lut_3_lut_4_lut_adj_299 (.A(n17458), .B(n17329), .C(n17327), 
         .D(n17273), .Z(n4311)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(570[10:40])
    defparam i1_2_lut_3_lut_4_lut_adj_299.init = 16'h2000;
    PFUMX i12487 (.BLUT(n16141), .ALUT(n16142), .C0(n17334), .Z(n16149));
    SPR16X4C Sprite_sizes_d12 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), .AD2(n17332), 
            .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4416), .DO0(n4410), 
            .DO1(n4411), .DO2(n4412), .DO3(n4413));
    defparam Sprite_sizes_d12.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d015 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4311), 
            .DO0(n4293), .DO1(n4294), .DO2(n4295), .DO3(n4296));
    defparam Sprite_positions_d015.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d014 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4311), 
            .DO0(n4297), .DO1(n4298), .DO2(n4299), .DO3(n4300));
    defparam Sprite_positions_d014.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d013 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4311), 
            .DO0(n4301), .DO1(n4302), .DO2(n4303), .DO3(n4304));
    defparam Sprite_positions_d013.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d012 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4276), 
            .DO0(n4258), .DO1(n4259), .DO2(n4260), .DO3(n4261));
    defparam Sprite_positions_d012.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d011 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4276), 
            .DO0(n4262), .DO1(n4263), .DO2(n4264), .DO3(n4265));
    defparam Sprite_positions_d011.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d010 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4276), 
            .DO0(n4266), .DO1(n4267), .DO2(n4268), .DO3(n4269));
    defparam Sprite_positions_d010.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d09 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4310), 
            .DO0(n4277), .DO1(n4278), .DO2(n4279), .DO3(n4280));
    defparam Sprite_positions_d09.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d08 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4310), 
            .DO0(n4281), .DO1(n4282), .DO2(n4283), .DO3(n4284));
    defparam Sprite_positions_d08.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d07 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), 
            .DI2(BUS_data[10]), .DI3(BUS_data[11]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4310), 
            .DO0(n4285), .DO1(n4286), .DO2(n4287), .DO3(n4288));
    defparam Sprite_positions_d07.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d06 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), 
            .DI2(BUS_data[2]), .DI3(BUS_data[3]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n3960), 
            .DO0(n4242), .DO1(n4243), .DO2(n4244), .DO3(n4245));
    defparam Sprite_positions_d06.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d05 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), 
            .DI2(BUS_data[6]), .DI3(BUS_data[7]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n3960), 
            .DO0(n4246), .DO1(n4247), .DO2(n4248), .DO3(n4249));
    defparam Sprite_positions_d05.initval = "0x0000000000000000";
    FADD2B mult_9u_9u_0_add_2_6 (.A0(s_mult_9u_9u_0_0_13), .A1(GND_net), 
           .B0(s_mult_9u_9u_0_1_13), .B1(s_mult_9u_9u_0_1_14), .CI(co_mult_9u_9u_0_2_5), 
           .COUT(co_mult_9u_9u_0_2_6), .S0(s_mult_9u_9u_0_2_13), .S1(s_mult_9u_9u_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 i7_4_lut (.A(currSprite[4]), .B(n14_adj_1917), .C(n15664), .D(currSprite[1]), 
         .Z(n70)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i7_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_rep_266_2_lut_4_lut (.A(n17314), .B(n17279), .C(n2539), 
         .D(n18260), .Z(n17274)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (B+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(458[95:155])
    defparam i1_2_lut_rep_266_2_lut_4_lut.init = 16'h3b00;
    PFUMX i12488 (.BLUT(n16143), .ALUT(n16144), .C0(n17334), .Z(n16150));
    SPR16X4C Sprite_positions_d00 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4310), 
            .DO0(n4289), .DO1(n4290), .DO2(n4291), .DO3(n4292));
    defparam Sprite_positions_d00.initval = "0x0000000000000000";
    LUT4 i12441_3_lut (.A(n4079), .B(n4095), .C(currSprite[4]), .Z(n16103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12441_3_lut.init = 16'hcaca;
    LUT4 i12440_3_lut (.A(n4044), .B(n4060), .C(currSprite[4]), .Z(n16102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12440_3_lut.init = 16'hcaca;
    PFUMX i12489 (.BLUT(n16145), .ALUT(n16146), .C0(n17334), .Z(n16151));
    SPR16X4C Sprite_positions_d03 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n3960), 
            .DO0(n4254), .DO1(n4255), .DO2(n4256), .DO3(n4257));
    defparam Sprite_positions_d03.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions_d01 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n17339), .AD1(n17333), 
            .AD2(n17332), .AD3(n17331), .CK(LOGIC_CLOCK), .WRE(n4276), 
            .DO0(n4270), .DO1(n4271), .DO2(n4272), .DO3(n4273));
    defparam Sprite_positions_d01.initval = "0x0000000000000000";
    DPR16X4C Sprite_options15 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4521), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4188));
    defparam Sprite_options15.initval = "0x0000000000000000";
    LUT4 i12431_3_lut (.A(n4076), .B(n4092), .C(currSprite[4]), .Z(n16093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12431_3_lut.init = 16'hcaca;
    DPR16X4C Sprite_options12 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4486), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4153));
    defparam Sprite_options12.initval = "0x0000000000000000";
    DPR16X4C Sprite_options9 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4520), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4172));
    defparam Sprite_options9.initval = "0x0000000000000000";
    LUT4 i12430_3_lut (.A(n4041), .B(n4057), .C(currSprite[4]), .Z(n16092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12430_3_lut.init = 16'hcaca;
    LUT4 i12428_3_lut (.A(n4075), .B(n4091), .C(currSprite[4]), .Z(n16090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12428_3_lut.init = 16'hcaca;
    DPR16X4C Sprite_options6 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4485), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4137));
    defparam Sprite_options6.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions3 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), 
            .WAD2(n17332), .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n3960), 
            .RAD0(currSprite[0]), .RAD1(currSprite[1]), .RAD2(currSprite[2]), 
            .RAD3(currSprite[3]), .DO0(n3939), .DO1(n3940), .DO2(n3941), 
            .DO3(n3942));
    defparam Sprite_positions3.initval = "0x0000000000000000";
    LUT4 i12427_3_lut (.A(n4040), .B(n4056), .C(currSprite[4]), .Z(n16089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12427_3_lut.init = 16'hcaca;
    PFUMX i12490 (.BLUT(n16147), .ALUT(n16148), .C0(n17334), .Z(n16152));
    CCU2D xPre_7__I_0_752_2 (.A0(xPre[0]), .B0(xOffset[0]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[1]), .B1(xOffset[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n14012), .S1(x[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(249[25:39])
    defparam xPre_7__I_0_752_2.INIT0 = 16'h7000;
    defparam xPre_7__I_0_752_2.INIT1 = 16'h5666;
    defparam xPre_7__I_0_752_2.INJECT1_0 = "NO";
    defparam xPre_7__I_0_752_2.INJECT1_1 = "NO";
    CCU2D add_617_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[0]), .B1(xOffset[0]), .C1(currColor[0]), .D1(GND_net), 
          .COUT(n14061), .S1(currAddress[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_1.INIT0 = 16'hF000;
    defparam add_617_1.INIT1 = 16'h9696;
    defparam add_617_1.INJECT1_0 = "NO";
    defparam add_617_1.INJECT1_1 = "NO";
    LUT4 i12418_3_lut (.A(n4074), .B(n4090), .C(currSprite[4]), .Z(n16080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12418_3_lut.init = 16'hcaca;
    LUT4 i12417_3_lut (.A(n4039), .B(n4055), .C(currSprite[4]), .Z(n16079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12417_3_lut.init = 16'hcaca;
    LUT4 LED_c_bdd_2_lut_3_lut (.A(n18256), .B(state[4]), .C(state[2]), 
         .Z(n18258)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam LED_c_bdd_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut (.A(currColor_lat[0]), .B(currColor_lat[1]), .C(currColor_lat[2]), 
         .D(currColor_lat[3]), .Z(n14447)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(359[9:29])
    defparam i1_3_lut_4_lut.init = 16'hfffb;
    LUT4 n15511_bdd_4_lut (.A(n17367), .B(n17275), .C(n17403), .D(n17405), 
         .Z(LOGIC_CLOCK_enable_33)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n15511_bdd_4_lut.init = 16'h0010;
    DPR16X4C Sprite_positions2 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), 
            .WAD2(n17332), .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4311), 
            .RAD0(currSprite[0]), .RAD1(currSprite[1]), .RAD2(currSprite[2]), 
            .RAD3(currSprite[3]), .DO0(n3990), .DO1(n3991), .DO2(n3992), 
            .DO3(n3993));
    defparam Sprite_positions2.initval = "0x0000000000000000";
    PFUMX i12502 (.BLUT(n16156), .ALUT(n16157), .C0(n17334), .Z(n16164));
    LUT4 i1_3_lut_4_lut_adj_300 (.A(currColor_lat[0]), .B(currColor_lat[1]), 
         .C(state[4]), .D(n15528), .Z(LOGIC_CLOCK_enable_140)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(359[9:29])
    defparam i1_3_lut_4_lut_adj_300.init = 16'h00f4;
    LUT4 i13060_4_lut (.A(n17306), .B(n16442), .C(Sprite_pointers_N_1136), 
         .D(n17287), .Z(LOGIC_CLOCK_enable_45)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i13060_4_lut.init = 16'h4000;
    FADD2B t_mult_9u_9u_0_add_3_5 (.A0(s_mult_9u_9u_0_2_15), .A1(s_mult_9u_9u_0_2_16), 
           .B0(mult_9u_9u_0_pp_4_15), .B1(mult_9u_9u_0_pp_4_16), .CI(co_t_mult_9u_9u_0_3_4), 
           .COUT(co_t_mult_9u_9u_0_3_5), .S0(RED_OUT_9__N_632[15]), .S1(RED_OUT_9__N_632[16])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 i12415_3_lut (.A(n4073), .B(n4089), .C(currSprite[4]), .Z(n16077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12415_3_lut.init = 16'hcaca;
    CCU2D add_10512_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14153), 
          .S0(n2539));
    defparam add_10512_cout.INIT0 = 16'h0000;
    defparam add_10512_cout.INIT1 = 16'h0000;
    defparam add_10512_cout.INJECT1_0 = "NO";
    defparam add_10512_cout.INJECT1_1 = "NO";
    LUT4 i12414_3_lut (.A(n4038), .B(n4054), .C(currSprite[4]), .Z(n16076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12414_3_lut.init = 16'hcaca;
    FADD2B mult_9u_9u_0_add_2_5 (.A0(s_mult_9u_9u_0_0_11), .A1(s_mult_9u_9u_0_0_12), 
           .B0(s_mult_9u_9u_0_1_11), .B1(s_mult_9u_9u_0_1_12), .CI(co_mult_9u_9u_0_2_4), 
           .COUT(co_mult_9u_9u_0_2_5), .S0(s_mult_9u_9u_0_2_11), .S1(s_mult_9u_9u_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_add_2_7_adj_301 (.A0(s_mult_10u_9u_0_0_15_adj_1920), 
           .A1(GND_net), .B0(s_mult_10u_9u_0_1_15_adj_1918), .B1(s_mult_10u_9u_0_1_16_adj_1919), 
           .CI(co_mult_10u_9u_0_2_6_adj_1914), .COUT(co_mult_10u_9u_0_2_7_adj_1921), 
           .S0(s_mult_10u_9u_0_2_15_adj_1922), .S1(s_mult_10u_9u_0_2_16_adj_1923)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_2_8_adj_302 (.A0(GND_net), .A1(GND_net), .B0(s_mult_10u_9u_0_1_17_adj_1924), 
           .B1(s_mult_10u_9u_0_1_18_adj_1925), .CI(co_mult_10u_9u_0_2_7_adj_1921), 
           .S0(s_mult_10u_9u_0_2_17_adj_1926), .S1(s_mult_10u_9u_0_2_18_adj_1927)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_1_7_adj_303 (.A0(GND_net), .A1(GND_net), .B0(mult_10u_9u_0_pp_3_17_adj_1929), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_1_6_adj_1928), .S0(s_mult_10u_9u_0_1_17_adj_1924), 
           .S1(s_mult_10u_9u_0_1_18_adj_1925)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_1_6_adj_304 (.A0(mult_10u_9u_0_pp_2_15_adj_1931), 
           .A1(GND_net), .B0(mult_10u_9u_0_pp_3_15_adj_1933), .B1(mult_10u_9u_0_pp_3_16_adj_1932), 
           .CI(co_mult_10u_9u_0_1_5_adj_1930), .COUT(co_mult_10u_9u_0_1_6_adj_1928), 
           .S0(s_mult_10u_9u_0_1_15_adj_1918), .S1(s_mult_10u_9u_0_1_16_adj_1919)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_1_5_adj_305 (.A0(mult_10u_9u_0_pp_2_13_adj_1936), 
           .A1(mult_10u_9u_0_pp_2_14_adj_1935), .B0(mult_10u_9u_0_pp_3_13_adj_1938), 
           .B1(mult_10u_9u_0_pp_3_14_adj_1937), .CI(co_mult_10u_9u_0_1_4_adj_1934), 
           .COUT(co_mult_10u_9u_0_1_5_adj_1930), .S0(s_mult_10u_9u_0_1_13_adj_1910), 
           .S1(s_mult_10u_9u_0_1_14_adj_1911)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_1_4_adj_306 (.A0(mult_10u_9u_0_pp_2_11_adj_1943), 
           .A1(mult_10u_9u_0_pp_2_12_adj_1942), .B0(mult_10u_9u_0_pp_3_11_adj_1945), 
           .B1(mult_10u_9u_0_pp_3_12_adj_1944), .CI(co_mult_10u_9u_0_1_3_adj_1939), 
           .COUT(co_mult_10u_9u_0_1_4_adj_1934), .S0(s_mult_10u_9u_0_1_11_adj_1940), 
           .S1(s_mult_10u_9u_0_1_12_adj_1941)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_1_3_adj_307 (.A0(mult_10u_9u_0_pp_2_9_adj_1950), 
           .A1(mult_10u_9u_0_pp_2_10_adj_1949), .B0(mult_10u_9u_0_pp_3_9_adj_1952), 
           .B1(mult_10u_9u_0_pp_3_10_adj_1951), .CI(co_mult_10u_9u_0_1_2_adj_1946), 
           .COUT(co_mult_10u_9u_0_1_3_adj_1939), .S0(s_mult_10u_9u_0_1_9_adj_1947), 
           .S1(s_mult_10u_9u_0_1_10_adj_1948)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_1_2_adj_308 (.A0(mult_10u_9u_0_pp_2_7_adj_1957), 
           .A1(mult_10u_9u_0_pp_2_8_adj_1956), .B0(mult_10u_9u_0_pp_3_7_adj_1959), 
           .B1(mult_10u_9u_0_pp_3_8_adj_1958), .CI(co_mult_10u_9u_0_1_1_adj_1953), 
           .COUT(co_mult_10u_9u_0_1_2_adj_1946), .S0(s_mult_10u_9u_0_1_7_adj_1954), 
           .S1(s_mult_10u_9u_0_1_8_adj_1955)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B Cadd_mult_10u_9u_0_1_1_adj_309 (.A0(GND_net), .A1(mult_10u_9u_0_pp_2_6_adj_1962), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_3_6_adj_1960), .CI(GND_net), 
           .COUT(co_mult_10u_9u_0_1_1_adj_1953), .S1(s_mult_10u_9u_0_1_6_adj_1961)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B Cadd_mult_10u_9u_0_0_8_adj_310 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_0_7_adj_1963), .S0(s_mult_10u_9u_0_0_15_adj_1920)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_0_7_adj_311 (.A0(GND_net), .A1(GND_net), .B0(mult_10u_9u_0_pp_1_13_adj_1965), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_0_6_adj_1964), .COUT(co_mult_10u_9u_0_0_7_adj_1963), 
           .S0(s_mult_10u_9u_0_0_13_adj_1912), .S1(s_mult_10u_9u_0_0_14_adj_1913)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    PFUMX i12503 (.BLUT(n16158), .ALUT(n16159), .C0(n17334), .Z(n16165));
    CCU2D sub_46_add_2_9 (.A0(currSprite_pos[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14060), .S0(SpriteRead_yInSprite[7]), .S1(SpriteRead_yValid_N_1156));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(272[44:107])
    defparam sub_46_add_2_9.INIT0 = 16'hf555;
    defparam sub_46_add_2_9.INIT1 = 16'h0000;
    defparam sub_46_add_2_9.INJECT1_0 = "NO";
    defparam sub_46_add_2_9.INJECT1_1 = "NO";
    FADD2B mult_9u_9u_0_add_2_4 (.A0(s_mult_9u_9u_0_0_9), .A1(s_mult_9u_9u_0_0_10), 
           .B0(s_mult_9u_9u_0_1_9), .B1(s_mult_9u_9u_0_1_10), .CI(co_mult_9u_9u_0_2_3), 
           .COUT(co_mult_9u_9u_0_2_4), .S0(s_mult_9u_9u_0_2_9), .S1(s_mult_9u_9u_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_add_0_6_adj_312 (.A0(mult_10u_9u_0_pp_0_11_adj_1967), 
           .A1(GND_net), .B0(mult_10u_9u_0_pp_1_11_adj_1971), .B1(mult_10u_9u_0_pp_1_12_adj_1970), 
           .CI(co_mult_10u_9u_0_0_5_adj_1966), .COUT(co_mult_10u_9u_0_0_6_adj_1964), 
           .S0(s_mult_10u_9u_0_0_11_adj_1968), .S1(s_mult_10u_9u_0_0_12_adj_1969)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    LUT4 i13059_4_lut (.A(n18260), .B(n14320), .C(n17428), .D(LOGIC_CLOCK_enable_52), 
         .Z(n16442)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i13059_4_lut.init = 16'h0004;
    FADD2B mult_10u_9u_0_add_0_5_adj_313 (.A0(mult_10u_9u_0_pp_0_9_adj_1976), 
           .A1(mult_10u_9u_0_pp_0_10_adj_1975), .B0(mult_10u_9u_0_pp_1_9_adj_1978), 
           .B1(mult_10u_9u_0_pp_1_10_adj_1977), .CI(co_mult_10u_9u_0_0_4_adj_1972), 
           .COUT(co_mult_10u_9u_0_0_5_adj_1966), .S0(s_mult_10u_9u_0_0_9_adj_1973), 
           .S1(s_mult_10u_9u_0_0_10_adj_1974)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    CCU2D add_19_2 (.A0(currSprite_pos[8]), .B0(currSprite_size[8]), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[9]), .B1(currSprite_size[9]), 
          .C1(GND_net), .D1(GND_net), .COUT(n14021), .S1(\SpriteRead_yValid_N_1158[1] ));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[132:154])
    defparam add_19_2.INIT0 = 16'h7000;
    defparam add_19_2.INIT1 = 16'h5666;
    defparam add_19_2.INJECT1_0 = "NO";
    defparam add_19_2.INJECT1_1 = "NO";
    FADD2B mult_9u_9u_0_add_1_6 (.A0(GND_net), .A1(GND_net), .B0(mult_9u_9u_0_pp_3_15), 
           .B1(mult_9u_9u_0_pp_3_16), .CI(co_mult_9u_9u_0_1_5), .COUT(co_mult_9u_9u_0_1_6), 
           .S0(s_mult_9u_9u_0_1_15), .S1(s_mult_9u_9u_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    LUT4 i12412_3_lut (.A(n4072), .B(n4088), .C(currSprite[4]), .Z(n16074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12412_3_lut.init = 16'hcaca;
    PFUMX i12504 (.BLUT(n16160), .ALUT(n16161), .C0(n17334), .Z(n16166));
    FD1P3DX ALPHA_WE_733 (.D(n18280), .SP(LOGIC_CLOCK_enable_45), .CK(LOGIC_CLOCK), 
            .CD(n17276), .Q(ALPHA_WE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam ALPHA_WE_733.GSR = "DISABLED";
    LUT4 i12411_3_lut (.A(n4037), .B(n4053), .C(currSprite[4]), .Z(n16073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12411_3_lut.init = 16'hcaca;
    PFUMX i12505 (.BLUT(n16162), .ALUT(n16163), .C0(n17334), .Z(n16167));
    LUT4 i12409_3_lut (.A(n4071), .B(n4087), .C(currSprite[4]), .Z(n16071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12409_3_lut.init = 16'hcaca;
    LUT4 i12408_3_lut (.A(n4036), .B(n4052), .C(currSprite[4]), .Z(n16070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12408_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut_then_4_lut (.A(n17382), .B(\BUS_ADDR_INTERNAL[3] ), 
         .C(\BUS_currGrantID[1] ), .D(\BUS_currGrantID[0] ), .Z(n17472)) /* synthesis lut_function=(A+!(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam i1_2_lut_rep_320_3_lut_4_lut_then_4_lut.init = 16'hafea;
    LUT4 i12406_3_lut (.A(n4070), .B(n4086), .C(currSprite[4]), .Z(n16068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12406_3_lut.init = 16'hcaca;
    LUT4 i12405_3_lut (.A(n4035), .B(n4051), .C(currSprite[4]), .Z(n16067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12405_3_lut.init = 16'hcaca;
    DPR16X4C Sprite_sizes15 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4416), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4083), .DO1(n4084), .DO2(n4085), .DO3(n4086));
    defparam Sprite_sizes15.initval = "0x0000000000000000";
    DPR16X4C Sprite_sizes14 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4416), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4087), .DO1(n4088), .DO2(n4089), .DO3(n4090));
    defparam Sprite_sizes14.initval = "0x0000000000000000";
    LUT4 i12403_3_lut (.A(n4069), .B(n4085), .C(currSprite[4]), .Z(n16065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12403_3_lut.init = 16'hcaca;
    CCU2D add_10512_13 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14152), .COUT(n14153));
    defparam add_10512_13.INIT0 = 16'heeee;
    defparam add_10512_13.INIT1 = 16'heeee;
    defparam add_10512_13.INJECT1_0 = "NO";
    defparam add_10512_13.INJECT1_1 = "NO";
    DPR16X4C Sprite_sizes13 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4416), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4091), .DO1(n4092), .DO2(n4093), .DO3(n4094));
    defparam Sprite_sizes13.initval = "0x0000000000000000";
    PFUMX i12517 (.BLUT(n16171), .ALUT(n16172), .C0(n17334), .Z(n16179));
    DPR16X4C Sprite_sizes12 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4381), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4048), .DO1(n4049), .DO2(n4050), .DO3(n4051));
    defparam Sprite_sizes12.initval = "0x0000000000000000";
    CCU2D add_10512_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[17]_adj_5 ), .D0(n18264), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), .D1(lastAddress_31__N_1310), 
          .CIN(n14151), .COUT(n14152));
    defparam add_10512_11.INIT0 = 16'h00ce;
    defparam add_10512_11.INIT1 = 16'hff20;
    defparam add_10512_11.INJECT1_0 = "NO";
    defparam add_10512_11.INJECT1_1 = "NO";
    FADD2B mult_10u_9u_0_add_0_4_adj_314 (.A0(mult_10u_9u_0_pp_0_7_adj_1983), 
           .A1(mult_10u_9u_0_pp_0_8_adj_1982), .B0(mult_10u_9u_0_pp_1_7_adj_1985), 
           .B1(mult_10u_9u_0_pp_1_8_adj_1984), .CI(co_mult_10u_9u_0_0_3_adj_1979), 
           .COUT(co_mult_10u_9u_0_0_4_adj_1972), .S0(s_mult_10u_9u_0_0_7_adj_1980), 
           .S1(s_mult_10u_9u_0_0_8_adj_1981)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    LUT4 i12402_3_lut (.A(n4034), .B(n4050), .C(currSprite[4]), .Z(n16064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12402_3_lut.init = 16'hcaca;
    DPR16X4C Sprite_sizes11 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4381), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4052), .DO1(n4053), .DO2(n4054), .DO3(n4055));
    defparam Sprite_sizes11.initval = "0x0000000000000000";
    CCU2D add_10512_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15]_adj_16 ), .D0(n18271), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16]_adj_15 ), 
          .D1(n18277), .CIN(n14150), .COUT(n14151));
    defparam add_10512_9.INIT0 = 16'hff31;
    defparam add_10512_9.INIT1 = 16'hff31;
    defparam add_10512_9.INJECT1_0 = "NO";
    defparam add_10512_9.INJECT1_1 = "NO";
    FADD2B mult_10u_9u_0_add_0_3_adj_315 (.A0(mult_10u_9u_0_pp_0_5_adj_1990), 
           .A1(mult_10u_9u_0_pp_0_6_adj_1989), .B0(mult_10u_9u_0_pp_1_5_adj_1992), 
           .B1(mult_10u_9u_0_pp_1_6_adj_1991), .CI(co_mult_10u_9u_0_0_2_adj_1986), 
           .COUT(co_mult_10u_9u_0_0_3_adj_1979), .S0(s_mult_10u_9u_0_0_5_adj_1987), 
           .S1(s_mult_10u_9u_0_0_6_adj_1988)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    CCU2D add_10512_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13]_adj_7 ), .D0(n18266), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14]_adj_3 ), 
          .D1(n18262), .CIN(n14149), .COUT(n14150));
    defparam add_10512_7.INIT0 = 16'h00ce;
    defparam add_10512_7.INIT1 = 16'h00ce;
    defparam add_10512_7.INJECT1_0 = "NO";
    defparam add_10512_7.INJECT1_1 = "NO";
    PFUMX i12518 (.BLUT(n16173), .ALUT(n16174), .C0(n17334), .Z(n16180));
    DPR16X4C Sprite_sizes10 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4381), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4056), .DO1(n4057), .DO2(n4058), .DO3(n4059));
    defparam Sprite_sizes10.initval = "0x0000000000000000";
    FADD2B mult_10u_9u_0_add_0_2_adj_316 (.A0(mult_10u_9u_0_pp_0_3_adj_1996), 
           .A1(mult_10u_9u_0_pp_0_4_adj_1995), .B0(mult_10u_9u_0_pp_1_3_adj_1998), 
           .B1(mult_10u_9u_0_pp_1_4_adj_1997), .CI(co_mult_10u_9u_0_0_1_adj_1993), 
           .COUT(co_mult_10u_9u_0_0_2_adj_1986), .S0(BLUE_OUT_9__N_687[3]), 
           .S1(s_mult_10u_9u_0_0_4_adj_1994)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    DPR16X4C Sprite_sizes9 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4415), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4067), .DO1(n4068), .DO2(n4069), .DO3(n4070));
    defparam Sprite_sizes9.initval = "0x0000000000000000";
    FADD2B Cadd_mult_10u_9u_0_0_1_adj_317 (.A0(GND_net), .A1(mult_10u_9u_0_pp_0_2_adj_2000), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_1_2_adj_1999), .CI(GND_net), 
           .COUT(co_mult_10u_9u_0_0_1_adj_1993), .S1(BLUE_OUT_9__N_687[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    DPR16X4C Sprite_sizes8 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4415), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4071), .DO1(n4072), .DO2(n4073), .DO3(n4074));
    defparam Sprite_sizes8.initval = "0x0000000000000000";
    FADD2B mult_10u_9u_0_Cadd_6_5_adj_318 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3_adj_2001), .S0(mult_10u_9u_0_pp_3_17_adj_1929)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    DPR16X4C Sprite_sizes7 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4415), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4075), .DO1(n4076), .DO2(n4077), .DO3(n4078));
    defparam Sprite_sizes7.initval = "0x0000000000000000";
    FADD2B mult_10u_9u_0_cin_lr_add_6_adj_319 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_6_adj_2002)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    DPR16X4C Sprite_sizes6 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4380), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4032), .DO1(n4033), .DO2(n4034), .DO3(n4035));
    defparam Sprite_sizes6.initval = "0x0000000000000000";
    FADD2B mult_10u_9u_0_Cadd_4_5_adj_320 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2_adj_2003), .S0(mult_10u_9u_0_pp_2_15_adj_1931)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    DPR16X4C Sprite_sizes5 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4380), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4036), .DO1(n4037), .DO2(n4038), .DO3(n4039));
    defparam Sprite_sizes5.initval = "0x0000000000000000";
    PFUMX i12519 (.BLUT(n16175), .ALUT(n16176), .C0(n17334), .Z(n16181));
    CCU2D add_10512_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n18273), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12]_adj_14 ), 
          .D1(n18272), .CIN(n14148), .COUT(n14149));
    defparam add_10512_5.INIT0 = 16'hff31;
    defparam add_10512_5.INIT1 = 16'h00ce;
    defparam add_10512_5.INJECT1_0 = "NO";
    defparam add_10512_5.INJECT1_1 = "NO";
    PFUMX i12520 (.BLUT(n16177), .ALUT(n16178), .C0(n17334), .Z(n16182));
    CCU2D add_10512_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[9]_adj_9 ), .D0(n18268), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n18269), 
          .CIN(n14147), .COUT(n14148));
    defparam add_10512_3.INIT0 = 16'h00ce;
    defparam add_10512_3.INIT1 = 16'h00ce;
    defparam add_10512_3.INJECT1_0 = "NO";
    defparam add_10512_3.INJECT1_1 = "NO";
    CCU2D add_10512_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8]_adj_8 ), 
          .D1(n18267), .COUT(n14147));
    defparam add_10512_1.INIT0 = 16'hF000;
    defparam add_10512_1.INIT1 = 16'h00ce;
    defparam add_10512_1.INJECT1_0 = "NO";
    defparam add_10512_1.INJECT1_1 = "NO";
    DPR16X4C Sprite_sizes0 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4415), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4079), .DO1(n4080), .DO2(n4081), .DO3(n4082));
    defparam Sprite_sizes0.initval = "0x0000000000000000";
    LUT4 inv_155_i1_1_lut_rep_431 (.A(xPre[0]), .Z(n17439)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i1_1_lut_rep_431.init = 16'h5555;
    PFUMX i12089 (.BLUT(n15749), .ALUT(n15750), .C0(n17334), .Z(Sprite_readData2_15__N_524[1]));
    LUT4 xPre_7__I_0_i4_4_lut_4_lut (.A(xPre[0]), .B(xPre[1]), .C(SpriteRead_xValid_N_1168[1]), 
         .D(SpriteRead_xValid_N_1168[0]), .Z(n4_c)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam xPre_7__I_0_i4_4_lut_4_lut.init = 16'h7130;
    PFUMX i12532 (.BLUT(n16186), .ALUT(n16187), .C0(n17334), .Z(n16194));
    PFUMX i12533 (.BLUT(n16188), .ALUT(n16189), .C0(n17334), .Z(n16195));
    PFUMX i12534 (.BLUT(n16190), .ALUT(n16191), .C0(n17334), .Z(n16196));
    LUT4 BUS_transferState_1__bdd_2_lut (.A(BUS_transferState[1]), .B(BUS_transferState[0]), 
         .Z(n16805)) /* synthesis lut_function=(A (B)) */ ;
    defparam BUS_transferState_1__bdd_2_lut.init = 16'h8888;
    DPR16X4C Sprite_sizes3 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4380), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4044), .DO1(n4045), .DO2(n4046), .DO3(n4047));
    defparam Sprite_sizes3.initval = "0x0000000000000000";
    DPR16X4C Sprite_sizes1 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4381), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4060), .DO1(n4061), .DO2(n4062), .DO3(n4063));
    defparam Sprite_sizes1.initval = "0x0000000000000000";
    LUT4 i11948_2_lut_rep_425_3_lut (.A(\state[0] ), .B(\state[1] ), .C(state[2]), 
         .Z(n17433)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i11948_2_lut_rep_425_3_lut.init = 16'h8080;
    DPR16X4C Sprite_sizes2 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4416), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n4095), .DO1(n4096), .DO2(n4097), .DO3(n4098));
    defparam Sprite_sizes2.initval = "0x0000000000000000";
    CCU2D xPre_7__I_0_752_6 (.A0(xPre[4]), .B0(xOffset_c[4]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[5]), .B1(xOffset_c[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14013), .COUT(n14014), .S0(x[4]), .S1(x[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(249[25:39])
    defparam xPre_7__I_0_752_6.INIT0 = 16'h5666;
    defparam xPre_7__I_0_752_6.INIT1 = 16'h5666;
    defparam xPre_7__I_0_752_6.INJECT1_0 = "NO";
    defparam xPre_7__I_0_752_6.INJECT1_1 = "NO";
    FD1P3DX BUS_transferState_i0 (.D(BUS_transferState_3__N_443[0]), .SP(LOGIC_CLOCK_enable_48), 
            .CK(LOGIC_CLOCK), .CD(n17276), .Q(BUS_transferState[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam BUS_transferState_i0.GSR = "DISABLED";
    CCU2D currSprite_999_add_4_9 (.A0(currSprite[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14133), .S0(n37[7]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999_add_4_9.INIT0 = 16'hfaaa;
    defparam currSprite_999_add_4_9.INIT1 = 16'h0000;
    defparam currSprite_999_add_4_9.INJECT1_0 = "NO";
    defparam currSprite_999_add_4_9.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_7 (.A0(SpriteRead_yInSprite_7__N_597[5]), .B0(currSprite_pos[13]), 
          .C0(GND_net), .D0(GND_net), .A1(SpriteRead_yInSprite_7__N_597[6]), 
          .B1(currSprite_pos[14]), .C1(GND_net), .D1(GND_net), .CIN(n14059), 
          .COUT(n14060), .S0(SpriteRead_yInSprite[5]), .S1(SpriteRead_yInSprite[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(272[44:107])
    defparam sub_46_add_2_7.INIT0 = 16'h5999;
    defparam sub_46_add_2_7.INIT1 = 16'h5999;
    defparam sub_46_add_2_7.INJECT1_0 = "NO";
    defparam sub_46_add_2_7.INJECT1_1 = "NO";
    FD1P3AX BUS_REQ_695 (.D(n14406), .SP(LOGIC_CLOCK_enable_49), .CK(LOGIC_CLOCK), 
            .Q(\BUS_currGrantID_3__N_74[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_REQ_695.GSR = "ENABLED";
    DPR16X4C Sprite_positions15 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4311), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3978), .DO1(n3979), .DO2(n3980), .DO3(n3981));
    defparam Sprite_positions15.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions14 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4311), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3982), .DO1(n3983), .DO2(n3984), .DO3(n3985));
    defparam Sprite_positions14.initval = "0x0000000000000000";
    CCU2D currSprite_999_add_4_7 (.A0(currSprite[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14132), .COUT(n14133), .S0(n37[5]), .S1(n37[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999_add_4_7.INIT0 = 16'hfaaa;
    defparam currSprite_999_add_4_7.INIT1 = 16'hfaaa;
    defparam currSprite_999_add_4_7.INJECT1_0 = "NO";
    defparam currSprite_999_add_4_7.INJECT1_1 = "NO";
    DPR16X4C Sprite_positions13 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4311), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3986), .DO1(n3987), .DO2(n3988), .DO3(n3989));
    defparam Sprite_positions13.initval = "0x0000000000000000";
    CCU2D sub_46_add_2_5 (.A0(MATRIX_CURRROW[3]), .B0(n17408), .C0(currSprite_pos[11]), 
          .D0(GND_net), .A1(MATRIX_CURRROW[4]), .B1(n17368), .C1(currSprite_pos[12]), 
          .D1(GND_net), .CIN(n14058), .COUT(n14059), .S0(SpriteRead_yInSprite[3]), 
          .S1(SpriteRead_yInSprite[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(272[44:107])
    defparam sub_46_add_2_5.INIT0 = 16'h9969;
    defparam sub_46_add_2_5.INIT1 = 16'h9969;
    defparam sub_46_add_2_5.INJECT1_0 = "NO";
    defparam sub_46_add_2_5.INJECT1_1 = "NO";
    LUT4 i2_2_lut_3_lut_3_lut_4_lut (.A(\state[0] ), .B(\state[1] ), .C(n17461), 
         .D(n17446), .Z(n6_adj_2004)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i2_2_lut_3_lut_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i1_2_lut_3_lut (.A(\state[0] ), .B(\state[1] ), .C(\state[3] ), 
         .Z(n6187)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    CCU2D currSprite_999_add_4_5 (.A0(currSprite[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14131), .COUT(n14132), .S0(n37[3]), .S1(n37[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999_add_4_5.INIT0 = 16'hfaaa;
    defparam currSprite_999_add_4_5.INIT1 = 16'hfaaa;
    defparam currSprite_999_add_4_5.INJECT1_0 = "NO";
    defparam currSprite_999_add_4_5.INJECT1_1 = "NO";
    DPR16X4C Sprite_positions12 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4276), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3943), .DO1(n3944), .DO2(n3945), .DO3(n3946));
    defparam Sprite_positions12.initval = "0x0000000000000000";
    LUT4 i2_2_lut_rep_380_3_lut_4_lut (.A(\state[0] ), .B(\state[1] ), .C(\state[3] ), 
         .D(state[2]), .Z(n17388)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_2_lut_rep_380_3_lut_4_lut.init = 16'h8000;
    PFUMX i12535 (.BLUT(n16192), .ALUT(n16193), .C0(n17334), .Z(n16197));
    LUT4 i6_1_lut_rep_434 (.A(\state[0] ), .Z(n17442)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i6_1_lut_rep_434.init = 16'h5555;
    CCU2D sub_46_add_2_3 (.A0(MATRIX_CURRROW[1]), .B0(MATRIX_CURRROW[0]), 
          .C0(currSprite_pos[9]), .D0(GND_net), .A1(MATRIX_CURRROW[2]), 
          .B1(n17452), .C1(currSprite_pos[10]), .D1(GND_net), .CIN(n14057), 
          .COUT(n14058), .S0(SpriteRead_yInSprite[1]), .S1(SpriteRead_yInSprite[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(272[44:107])
    defparam sub_46_add_2_3.INIT0 = 16'h9969;
    defparam sub_46_add_2_3.INIT1 = 16'h9969;
    defparam sub_46_add_2_3.INJECT1_0 = "NO";
    defparam sub_46_add_2_3.INJECT1_1 = "NO";
    FD1P3AX frameEndClock_700 (.D(n18280), .SP(LOGIC_CLOCK_enable_50), .CK(LOGIC_CLOCK), 
            .Q(frameEndClock)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam frameEndClock_700.GSR = "ENABLED";
    DPR16X4C Sprite_positions11 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4276), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3947), .DO1(n3948), .DO2(n3949), .DO3(n3950));
    defparam Sprite_positions11.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions10 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4276), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3951), .DO1(n3952), .DO2(n3953), .DO3(n3954));
    defparam Sprite_positions10.initval = "0x0000000000000000";
    CCU2D currSprite_999_add_4_3 (.A0(currSprite[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14130), .COUT(n14131), .S0(n37[1]), .S1(n37[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999_add_4_3.INIT0 = 16'hfaaa;
    defparam currSprite_999_add_4_3.INIT1 = 16'hfaaa;
    defparam currSprite_999_add_4_3.INJECT1_0 = "NO";
    defparam currSprite_999_add_4_3.INJECT1_1 = "NO";
    CCU2D sub_46_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(MATRIX_CURRROW[0]), .B1(currSprite_pos[8]), .C1(GND_net), 
          .D1(GND_net), .COUT(n14057), .S1(SpriteRead_yInSprite[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(272[44:107])
    defparam sub_46_add_2_1.INIT0 = 16'h0000;
    defparam sub_46_add_2_1.INIT1 = 16'ha666;
    defparam sub_46_add_2_1.INJECT1_0 = "NO";
    defparam sub_46_add_2_1.INJECT1_1 = "NO";
    CCU2D BLUE_OUT_9__I_0_20 (.A0(BLUE_OUT_9__N_687[18]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14056), .S0(BLUE_OUT[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_20.INIT0 = 16'h5aaa;
    defparam BLUE_OUT_9__I_0_20.INIT1 = 16'h0000;
    defparam BLUE_OUT_9__I_0_20.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_20.INJECT1_1 = "NO";
    DPR16X4C Sprite_positions9 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4310), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3962), .DO1(n3963), .DO2(n3964), .DO3(n3965));
    defparam Sprite_positions9.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions8 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4310), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3966), .DO1(n3967), .DO2(n3968), .DO3(n3969));
    defparam Sprite_positions8.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions7 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4310), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3970), .DO1(n3971), .DO2(n3972), .DO3(n3973));
    defparam Sprite_positions7.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions6 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n3960), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3927), .DO1(n3928), .DO2(n3929), .DO3(n3930));
    defparam Sprite_positions6.initval = "0x0000000000000000";
    DPR16X4C Sprite_positions5 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .WAD0(n17339), .WAD1(n17333), .WAD2(n17332), 
            .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n3960), .RAD0(currSprite[0]), 
            .RAD1(currSprite[1]), .RAD2(currSprite[2]), .RAD3(currSprite[3]), 
            .DO0(n3931), .DO1(n3932), .DO2(n3933), .DO3(n3934));
    defparam Sprite_positions5.initval = "0x0000000000000000";
    LUT4 i6_4_lut (.A(currSprite[6]), .B(currSprite[7]), .C(currSprite[3]), 
         .D(currSprite[5]), .Z(n14_adj_1917)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i6_4_lut.init = 16'hfeff;
    PFUMX i12547 (.BLUT(n16201), .ALUT(n16202), .C0(n17334), .Z(n16209));
    LUT4 i1_4_lut_4_lut (.A(\state[0] ), .B(n17451), .C(n17468), .D(state[4]), 
         .Z(n60_adj_2005)) /* synthesis lut_function=(A (B (C (D)))+!A (D)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_4_lut.init = 16'hd500;
    LUT4 i1_2_lut_4_lut_4_lut (.A(\state[0] ), .B(state[4]), .C(n17429), 
         .D(n15442), .Z(LOGIC_CLOCK_enable_38)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 state_7__I_0_770_i13_2_lut_rep_435 (.A(state[6]), .B(state[7]), 
         .Z(n17443)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(381[10:23])
    defparam state_7__I_0_770_i13_2_lut_rep_435.init = 16'hbbbb;
    PFUMX i12548 (.BLUT(n16203), .ALUT(n16204), .C0(n17334), .Z(n16210));
    LUT4 i12400_3_lut (.A(n4068), .B(n4084), .C(currSprite[4]), .Z(n16062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12400_3_lut.init = 16'hcaca;
    LUT4 i12004_2_lut (.A(currSprite[0]), .B(currSprite[2]), .Z(n15664)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12004_2_lut.init = 16'h8888;
    DPR16X4C Sprite_positions0 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .WAD0(n17339), .WAD1(n17333), 
            .WAD2(n17332), .WAD3(n17331), .WCK(LOGIC_CLOCK), .WRE(n4310), 
            .RAD0(currSprite[0]), .RAD1(currSprite[1]), .RAD2(currSprite[2]), 
            .RAD3(currSprite[3]), .DO0(n3974), .DO1(n3975), .DO2(n3976), 
            .DO3(n3977));
    defparam Sprite_positions0.initval = "0x0000000000000000";
    CCU2D currSprite_999_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n14130), .S1(n37[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999_add_4_1.INIT0 = 16'hF000;
    defparam currSprite_999_add_4_1.INIT1 = 16'h0555;
    defparam currSprite_999_add_4_1.INJECT1_0 = "NO";
    defparam currSprite_999_add_4_1.INJECT1_1 = "NO";
    PFUMX i12549 (.BLUT(n16205), .ALUT(n16206), .C0(n17334), .Z(n16211));
    LUT4 i12399_3_lut (.A(n4033), .B(n4049), .C(currSprite[4]), .Z(n16061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12399_3_lut.init = 16'hcaca;
    LUT4 i12394_3_lut (.A(n4082), .B(n4098), .C(currSprite[4]), .Z(n16056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12394_3_lut.init = 16'hcaca;
    LUT4 i12393_3_lut (.A(n4047), .B(n4063), .C(currSprite[4]), .Z(n16055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12393_3_lut.init = 16'hcaca;
    LUT4 i12391_3_lut (.A(n4172), .B(n4188), .C(currSprite[4]), .Z(n16053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12391_3_lut.init = 16'hcaca;
    PFUMX i12550 (.BLUT(n16207), .ALUT(n16208), .C0(n17334), .Z(n16212));
    LUT4 i12390_3_lut (.A(n4137), .B(n4153), .C(currSprite[4]), .Z(n16052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12390_3_lut.init = 16'hcaca;
    LUT4 i13106_3_lut_rep_268_4_lut (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), 
         .B(n2504), .C(n2539), .D(n17314), .Z(n17276)) /* synthesis lut_function=(A (B (C+!(D)))+!A (C+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(458[95:155])
    defparam i13106_3_lut_rep_268_4_lut.init = 16'hd0dd;
    FADD2B mult_10u_9u_0_cin_lr_add_4_adj_321 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_4_adj_2006)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_Cadd_2_5_adj_322 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1_adj_2007), .S0(mult_10u_9u_0_pp_1_13_adj_1965)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_cin_lr_add_2_adj_323 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_2_adj_2008)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_Cadd_0_5_adj_324 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_adj_2009), .S0(mult_10u_9u_0_pp_0_11_adj_1967)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    PFUMX i12092 (.BLUT(n15752), .ALUT(n15753), .C0(n17334), .Z(Sprite_readData2_15__N_524[2]));
    LUT4 i1_2_lut_4_lut (.A(n17374), .B(n17458), .C(n17373), .D(Sprite_pointers_N_1123), 
         .Z(n4626)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A !(B+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(573[21:66])
    defparam i1_2_lut_4_lut.init = 16'hb300;
    LUT4 i12388_3_lut (.A(n4077), .B(n4093), .C(currSprite[4]), .Z(n16050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12388_3_lut.init = 16'hcaca;
    FADD2B mult_9u_9u_0_add_2_3 (.A0(s_mult_9u_9u_0_0_7), .A1(s_mult_9u_9u_0_0_8), 
           .B0(s_mult_9u_9u_0_1_7), .B1(s_mult_9u_9u_0_1_8), .CI(co_mult_9u_9u_0_2_2), 
           .COUT(co_mult_9u_9u_0_2_3), .S0(RED_OUT_9__N_632[7]), .S1(s_mult_9u_9u_0_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    AND2 AND2_t13_adj_325 (.A(VRAM_DATA_OUT[20]), .B(RED_OUT_9__N_768[0]), 
         .Z(BLUE_OUT_9__N_687[0])) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(170[10:65])
    AND2 AND2_t12_adj_326 (.A(VRAM_DATA_OUT[20]), .B(RED_OUT_9__N_768[2]), 
         .Z(mult_10u_9u_0_pp_1_2_adj_1999)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(172[10:65])
    AND2 AND2_t11_adj_327 (.A(VRAM_DATA_OUT[20]), .B(RED_OUT_9__N_768[4]), 
         .Z(mult_10u_9u_0_pp_2_4_adj_2010)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(174[10:65])
    AND2 AND2_t10_adj_328 (.A(VRAM_DATA_OUT[20]), .B(RED_OUT_9__N_768[6]), 
         .Z(mult_10u_9u_0_pp_3_6_adj_1960)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(176[10:65])
    FADD2B mult_9u_9u_0_cin_lr_add_0_adj_329 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_0_adj_2011)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    AND2 AND2_t0_adj_330 (.A(GREEN_READ[8]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_16_adj_2012)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(183[10:64])
    AND2 AND2_t1_adj_331 (.A(GREEN_READ[7]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_15_adj_2013)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(181[10:64])
    AND2 AND2_t2_adj_332 (.A(GREEN_READ[6]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_14_adj_2014)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(179[10:64])
    FD1P3AX SpriteLut_writeClk_741 (.D(Sprite_writeClk_N_1144), .SP(LOGIC_CLOCK_enable_51), 
            .CK(LOGIC_CLOCK), .Q(SpriteLut_writeClk)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam SpriteLut_writeClk_741.GSR = "DISABLED";
    FD1P3DX GR_WR_CLK_728 (.D(GR_WR_CLK_N_1081), .SP(LOGIC_CLOCK_enable_52), 
            .CK(LOGIC_CLOCK), .CD(n17276), .Q(GR_WR_CLK)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_CLK_728.GSR = "DISABLED";
    FD1P3DX GREEN_WE_731 (.D(n18280), .SP(LOGIC_CLOCK_enable_53), .CK(LOGIC_CLOCK), 
            .CD(n17276), .Q(GREEN_WE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GREEN_WE_731.GSR = "DISABLED";
    FD1P3DX BLUE_WE_732 (.D(n18280), .SP(LOGIC_CLOCK_enable_54), .CK(LOGIC_CLOCK), 
            .CD(n17276), .Q(BLUE_WE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam BLUE_WE_732.GSR = "DISABLED";
    LUT4 i10543_3_lut_4_lut (.A(currColor[1]), .B(currColor[0]), .C(currColor[2]), 
         .D(currColor[3]), .Z(n3[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10543_3_lut_4_lut.init = 16'h7f80;
    CCU2D add_1840_9 (.A0(x[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14129), 
          .S0(currAddress_17__N_742[8]), .S1(currAddress_17__N_742[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[150:167])
    defparam add_1840_9.INIT0 = 16'h5aaa;
    defparam add_1840_9.INIT1 = 16'h0000;
    defparam add_1840_9.INJECT1_0 = "NO";
    defparam add_1840_9.INJECT1_1 = "NO";
    AND2 AND2_t3_adj_333 (.A(GREEN_READ[5]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_13_adj_2015)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(177[10:64])
    CCU2D BLUE_OUT_9__I_0_18 (.A0(BLUE_OUT_9__N_687[16]), .B0(BLUE_OUT_9__N_706[16]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[17]), .B1(BLUE_OUT_9__N_706[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14055), .COUT(n14056), .S0(BLUE_OUT[7]), 
          .S1(BLUE_OUT[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_18.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_18.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_18.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_18.INJECT1_1 = "NO";
    AND2 AND2_t4_adj_334 (.A(GREEN_READ[4]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_12_adj_2016)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(175[10:64])
    AND2 AND2_t5_adj_335 (.A(GREEN_READ[3]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_11_adj_2017)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(173[10:64])
    AND2 AND2_t6_adj_336 (.A(GREEN_READ[2]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_10_adj_2018)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(171[10:64])
    CCU2D yPre_7__I_0_757_9 (.A0(yOffset_c[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14019), .S0(y[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[24:38])
    defparam yPre_7__I_0_757_9.INIT0 = 16'hfaaa;
    defparam yPre_7__I_0_757_9.INIT1 = 16'h0000;
    defparam yPre_7__I_0_757_9.INJECT1_0 = "NO";
    defparam yPre_7__I_0_757_9.INJECT1_1 = "NO";
    LUT4 i10536_2_lut_3_lut (.A(currColor[1]), .B(currColor[0]), .C(currColor[2]), 
         .Z(n3[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10536_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_4_lut_4_lut_adj_337 (.A(state[4]), .B(n73), .C(n17402), .D(n17406), 
         .Z(n62)) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i1_4_lut_4_lut_adj_337.init = 16'hf444;
    AND2 AND2_t7_adj_338 (.A(GREEN_READ[1]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_9_adj_2019)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(169[10:63])
    MULT2 mult_9u_9u_0_mult_6_4_adj_339 (.A0(GREEN_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), 
          .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), .CI(mco_15_adj_2022), 
          .P0(mult_9u_9u_0_pp_3_15_adj_2021), .P1(mult_9u_9u_0_pp_3_16_adj_2020)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 SRAM_WE_N_1255_I_0_301_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17371), .D(n18270), .Z(lastAddress_31__N_1425)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_301_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 i2_4_lut_4_lut_4_lut (.A(state[4]), .B(\state[1] ), .C(n8405), 
         .D(\state[0] ), .Z(n14339)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i2_4_lut_4_lut_4_lut.init = 16'h4044;
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[4]), .B(n17403), .C(n17447), .D(state[5]), 
         .Z(n15_adj_2023)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hfffd;
    MULT2 mult_9u_9u_0_mult_6_3_adj_340 (.A0(GREEN_READ[6]), .A1(GREEN_READ[7]), 
          .A2(GREEN_READ[7]), .A3(GREEN_READ[8]), .B0(ALPHA_READ[7]), 
          .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), 
          .CI(mco_14_adj_2026), .CO(mco_15_adj_2022), .P0(mult_9u_9u_0_pp_3_13_adj_2025), 
          .P1(mult_9u_9u_0_pp_3_14_adj_2024)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 i1_2_lut_3_lut_4_lut_adj_341 (.A(n17385), .B(n17384), .C(n6250), 
         .D(n17458), .Z(LOGIC_CLOCK_enable_74)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(570[10:40])
    defparam i1_2_lut_3_lut_4_lut_adj_341.init = 16'h1000;
    LUT4 i1_2_lut_rep_303_3_lut_4_lut (.A(n17385), .B(n17384), .C(n17382), 
         .D(n17371), .Z(n17311)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(570[10:40])
    defparam i1_2_lut_rep_303_3_lut_4_lut.init = 16'hfffe;
    FD1P3AX GR_WR_DOUT_16__i10 (.D(GR_WR_DOUT[9]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i10.GSR = "DISABLED";
    FD1P3AX GR_WR_DOUT_16__i9 (.D(GR_WR_DOUT[8]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i9.GSR = "DISABLED";
    MULT2 mult_9u_9u_0_mult_6_2_adj_342 (.A0(GREEN_READ[4]), .A1(GREEN_READ[5]), 
          .A2(GREEN_READ[5]), .A3(GREEN_READ[6]), .B0(ALPHA_READ[7]), 
          .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), 
          .CI(mco_13_adj_2029), .CO(mco_14_adj_2026), .P0(mult_9u_9u_0_pp_3_11_adj_2028), 
          .P1(mult_9u_9u_0_pp_3_12_adj_2027)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_6_1_adj_343 (.A0(GREEN_READ[2]), .A1(GREEN_READ[3]), 
          .A2(GREEN_READ[3]), .A3(GREEN_READ[4]), .B0(ALPHA_READ[7]), 
          .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), 
          .CI(mco_12_adj_2032), .CO(mco_13_adj_2029), .P0(mult_9u_9u_0_pp_3_9_adj_2031), 
          .P1(mult_9u_9u_0_pp_3_10_adj_2030)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_6_0_adj_344 (.A0(GREEN_READ[0]), .A1(GREEN_READ[1]), 
          .A2(GREEN_READ[1]), .A3(GREEN_READ[2]), .B0(ALPHA_READ[7]), 
          .B1(ALPHA_READ[6]), .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), 
          .CI(mult_9u_9u_0_cin_lr_6_adj_2035), .CO(mco_12_adj_2032), .P0(mult_9u_9u_0_pp_3_7_adj_2034), 
          .P1(mult_9u_9u_0_pp_3_8_adj_2033)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FD1P3AX GR_WR_DOUT_16__i8 (.D(GR_WR_DOUT[7]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i8.GSR = "DISABLED";
    MULT2 mult_9u_9u_0_mult_4_4_adj_345 (.A0(GREEN_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), 
          .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), .CI(mco_11_adj_2038), 
          .P0(mult_9u_9u_0_pp_2_13_adj_2037), .P1(mult_9u_9u_0_pp_2_14_adj_2036)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FD1P3AX GR_WR_DOUT_16__i7 (.D(GR_WR_DOUT[6]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i7.GSR = "DISABLED";
    PFUMX i12095 (.BLUT(n15755), .ALUT(n15756), .C0(n17334), .Z(Sprite_readData2_15__N_524[3]));
    LUT4 i12387_3_lut (.A(n4042), .B(n4058), .C(currSprite[4]), .Z(n16049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12387_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut_4_lut (.A(state[4]), .B(state[6]), .C(state[7]), .D(\state[3] ), 
         .Z(n10)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i4_4_lut_4_lut.init = 16'hf7ff;
    MULT2 mult_9u_9u_0_mult_4_3_adj_346 (.A0(GREEN_READ[6]), .A1(GREEN_READ[7]), 
          .A2(GREEN_READ[7]), .A3(GREEN_READ[8]), .B0(ALPHA_READ[5]), 
          .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), 
          .CI(mco_10_adj_2041), .CO(mco_11_adj_2038), .P0(mult_9u_9u_0_pp_2_11_adj_2040), 
          .P1(mult_9u_9u_0_pp_2_12_adj_2039)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B t_mult_9u_9u_0_add_3_4 (.A0(s_mult_9u_9u_0_2_13), .A1(s_mult_9u_9u_0_2_14), 
           .B0(mult_9u_9u_0_pp_4_13), .B1(mult_9u_9u_0_pp_4_14), .CI(co_t_mult_9u_9u_0_3_3), 
           .COUT(co_t_mult_9u_9u_0_3_4), .S0(RED_OUT_9__N_632[13]), .S1(RED_OUT_9__N_632[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_4_2_adj_347 (.A0(GREEN_READ[4]), .A1(GREEN_READ[5]), 
          .A2(GREEN_READ[5]), .A3(GREEN_READ[6]), .B0(ALPHA_READ[5]), 
          .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), 
          .CI(mco_9_adj_2044), .CO(mco_10_adj_2041), .P0(mult_9u_9u_0_pp_2_9_adj_2043), 
          .P1(mult_9u_9u_0_pp_2_10_adj_2042)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 i12385_3_lut (.A(n3972), .B(n3988), .C(currSprite[4]), .Z(n16047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12385_3_lut.init = 16'hcaca;
    CCU2D add_1840_7 (.A0(x[5]), .B0(x[6]), .C0(GND_net), .D0(GND_net), 
          .A1(x[6]), .B1(x[7]), .C1(GND_net), .D1(GND_net), .CIN(n14128), 
          .COUT(n14129), .S0(currAddress_17__N_742[6]), .S1(currAddress_17__N_742[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[150:167])
    defparam add_1840_7.INIT0 = 16'h5666;
    defparam add_1840_7.INIT1 = 16'h5666;
    defparam add_1840_7.INJECT1_0 = "NO";
    defparam add_1840_7.INJECT1_1 = "NO";
    CCU2D BLUE_OUT_9__I_0_16 (.A0(BLUE_OUT_9__N_687[14]), .B0(BLUE_OUT_9__N_706[14]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[15]), .B1(BLUE_OUT_9__N_706[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14054), .COUT(n14055), .S0(BLUE_OUT[5]), 
          .S1(BLUE_OUT[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_16.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_16.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_16.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_16.INJECT1_1 = "NO";
    CCU2D yPre_7__I_0_757_7 (.A0(yOffset_c[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(yOffset_c[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14018), .COUT(n14019), .S0(y[5]), .S1(y[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[24:38])
    defparam yPre_7__I_0_757_7.INIT0 = 16'hfaaa;
    defparam yPre_7__I_0_757_7.INIT1 = 16'hfaaa;
    defparam yPre_7__I_0_757_7.INJECT1_0 = "NO";
    defparam yPre_7__I_0_757_7.INJECT1_1 = "NO";
    CCU2D yPre_7__I_0_757_5 (.A0(MATRIX_CURRROW[3]), .B0(n17408), .C0(\yOffset[3] ), 
          .D0(GND_net), .A1(MATRIX_CURRROW[4]), .B1(n17368), .C1(yOffset_c[4]), 
          .D1(GND_net), .CIN(n14017), .COUT(n14018), .S0(y[3]), .S1(y[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[24:38])
    defparam yPre_7__I_0_757_5.INIT0 = 16'h9696;
    defparam yPre_7__I_0_757_5.INIT1 = 16'h9696;
    defparam yPre_7__I_0_757_5.INJECT1_0 = "NO";
    defparam yPre_7__I_0_757_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_348 (.A(n17458), .B(n17329), .C(n17312), .D(n6250), 
         .Z(LOGIC_CLOCK_enable_53)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(570[10:40])
    defparam i2_3_lut_4_lut_adj_348.init = 16'h0d00;
    MULT2 mult_9u_9u_0_mult_4_1_adj_349 (.A0(GREEN_READ[2]), .A1(GREEN_READ[3]), 
          .A2(GREEN_READ[3]), .A3(GREEN_READ[4]), .B0(ALPHA_READ[5]), 
          .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), 
          .CI(mco_8_adj_2047), .CO(mco_9_adj_2044), .P0(mult_9u_9u_0_pp_2_7_adj_2046), 
          .P1(mult_9u_9u_0_pp_2_8_adj_2045)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_4_0_adj_350 (.A0(GREEN_READ[0]), .A1(GREEN_READ[1]), 
          .A2(GREEN_READ[1]), .A3(GREEN_READ[2]), .B0(ALPHA_READ[5]), 
          .B1(ALPHA_READ[4]), .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), 
          .CI(mult_9u_9u_0_cin_lr_4_adj_2050), .CO(mco_8_adj_2047), .P0(mult_9u_9u_0_pp_2_5_adj_2049), 
          .P1(mult_9u_9u_0_pp_2_6_adj_2048)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_2_4_adj_351 (.A0(GREEN_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), 
          .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), .CI(mco_7_adj_2053), 
          .P0(mult_9u_9u_0_pp_1_11_adj_2052), .P1(mult_9u_9u_0_pp_1_12_adj_2051)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_2_3_adj_352 (.A0(GREEN_READ[6]), .A1(GREEN_READ[7]), 
          .A2(GREEN_READ[7]), .A3(GREEN_READ[8]), .B0(ALPHA_READ[3]), 
          .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), 
          .CI(mco_6_adj_2056), .CO(mco_7_adj_2053), .P0(mult_9u_9u_0_pp_1_9_adj_2055), 
          .P1(mult_9u_9u_0_pp_1_10_adj_2054)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_2_2_adj_353 (.A0(GREEN_READ[4]), .A1(GREEN_READ[5]), 
          .A2(GREEN_READ[5]), .A3(GREEN_READ[6]), .B0(ALPHA_READ[3]), 
          .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), 
          .CI(mco_5_adj_2059), .CO(mco_6_adj_2056), .P0(mult_9u_9u_0_pp_1_7_adj_2058), 
          .P1(mult_9u_9u_0_pp_1_8_adj_2057)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B t_mult_9u_9u_0_add_3_3 (.A0(s_mult_9u_9u_0_2_11), .A1(s_mult_9u_9u_0_2_12), 
           .B0(mult_9u_9u_0_pp_4_11), .B1(mult_9u_9u_0_pp_4_12), .CI(co_t_mult_9u_9u_0_3_2), 
           .COUT(co_t_mult_9u_9u_0_3_3), .S0(RED_OUT_9__N_632[11]), .S1(RED_OUT_9__N_632[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_9u_9u_0_mult_2_1_adj_354 (.A0(GREEN_READ[2]), .A1(GREEN_READ[3]), 
          .A2(GREEN_READ[3]), .A3(GREEN_READ[4]), .B0(ALPHA_READ[3]), 
          .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), 
          .CI(mco_4_adj_2062), .CO(mco_5_adj_2059), .P0(mult_9u_9u_0_pp_1_5_adj_2061), 
          .P1(mult_9u_9u_0_pp_1_6_adj_2060)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 i13029_4_lut_4_lut (.A(state[4]), .B(n15378), .C(n95), .D(n17349), 
         .Z(state_7__N_336[4])) /* synthesis lut_function=(!(A (C (D))+!A (B (D)+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i13029_4_lut_4_lut.init = 16'h0bff;
    LUT4 i12384_3_lut (.A(n3937), .B(n3953), .C(currSprite[4]), .Z(n16046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12384_3_lut.init = 16'hcaca;
    LUT4 i12382_3_lut (.A(n3977), .B(n3993), .C(currSprite[4]), .Z(n16044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12382_3_lut.init = 16'hcaca;
    LUT4 i12381_3_lut (.A(n3942), .B(n3958), .C(currSprite[4]), .Z(n16043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12381_3_lut.init = 16'hcaca;
    MULT2 mult_9u_9u_0_mult_2_0_adj_355 (.A0(GREEN_READ[0]), .A1(GREEN_READ[1]), 
          .A2(GREEN_READ[1]), .A3(GREEN_READ[2]), .B0(ALPHA_READ[3]), 
          .B1(ALPHA_READ[2]), .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), 
          .CI(mult_9u_9u_0_cin_lr_2_adj_2065), .CO(mco_4_adj_2062), .P0(mult_9u_9u_0_pp_1_3_adj_2064), 
          .P1(mult_9u_9u_0_pp_1_4_adj_2063)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_0_4_adj_356 (.A0(GREEN_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), 
          .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), .CI(mco_3_adj_2068), 
          .P0(mult_9u_9u_0_pp_0_9_adj_2067), .P1(mult_9u_9u_0_pp_0_10_adj_2066)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    CCU2D add_1840_5 (.A0(x[3]), .B0(x[4]), .C0(GND_net), .D0(GND_net), 
          .A1(x[4]), .B1(x[5]), .C1(GND_net), .D1(GND_net), .CIN(n14127), 
          .COUT(n14128), .S0(currAddress_17__N_742[4]), .S1(currAddress_17__N_742[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[150:167])
    defparam add_1840_5.INIT0 = 16'h5666;
    defparam add_1840_5.INIT1 = 16'h5666;
    defparam add_1840_5.INJECT1_0 = "NO";
    defparam add_1840_5.INJECT1_1 = "NO";
    FD1P3DX RED_WE_730 (.D(n18280), .SP(LOGIC_CLOCK_enable_74), .CK(LOGIC_CLOCK), 
            .CD(n17276), .Q(RED_WE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam RED_WE_730.GSR = "DISABLED";
    MULT2 mult_9u_9u_0_mult_0_3_adj_357 (.A0(GREEN_READ[6]), .A1(GREEN_READ[7]), 
          .A2(GREEN_READ[7]), .A3(GREEN_READ[8]), .B0(ALPHA_READ[1]), 
          .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), 
          .CI(mco_2_adj_2071), .CO(mco_3_adj_2068), .P0(mult_9u_9u_0_pp_0_7_adj_2070), 
          .P1(mult_9u_9u_0_pp_0_8_adj_2069)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 state_7__I_0_771_i12_2_lut_rep_389_2_lut (.A(state[4]), .B(state[5]), 
         .Z(n17397)) /* synthesis lut_function=((B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam state_7__I_0_771_i12_2_lut_rep_389_2_lut.init = 16'hdddd;
    CCU2D BLUE_OUT_9__I_0_14 (.A0(BLUE_OUT_9__N_687[12]), .B0(BLUE_OUT_9__N_706[12]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[13]), .B1(BLUE_OUT_9__N_706[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14053), .COUT(n14054), .S0(BLUE_OUT[3]), 
          .S1(BLUE_OUT[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_14.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_14.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_14.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_14.INJECT1_1 = "NO";
    PFUMX i12098 (.BLUT(n15758), .ALUT(n15759), .C0(n17334), .Z(Sprite_readData2_15__N_524[4]));
    MULT2 mult_9u_9u_0_mult_0_2_adj_358 (.A0(GREEN_READ[4]), .A1(GREEN_READ[5]), 
          .A2(GREEN_READ[5]), .A3(GREEN_READ[6]), .B0(ALPHA_READ[1]), 
          .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), 
          .CI(mco_1_adj_2074), .CO(mco_2_adj_2071), .P0(mult_9u_9u_0_pp_0_5_adj_2073), 
          .P1(mult_9u_9u_0_pp_0_6_adj_2072)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    CCU2D yPre_7__I_0_757_3 (.A0(MATRIX_CURRROW[1]), .B0(MATRIX_CURRROW[0]), 
          .C0(\yOffset[1] ), .D0(GND_net), .A1(MATRIX_CURRROW[2]), .B1(n17452), 
          .C1(\yOffset[2] ), .D1(GND_net), .CIN(n14016), .COUT(n14017), 
          .S0(y[1]), .S1(y[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[24:38])
    defparam yPre_7__I_0_757_3.INIT0 = 16'h9696;
    defparam yPre_7__I_0_757_3.INIT1 = 16'h9696;
    defparam yPre_7__I_0_757_3.INJECT1_0 = "NO";
    defparam yPre_7__I_0_757_3.INJECT1_1 = "NO";
    FD1P3AX GR_WR_DOUT_16__i6 (.D(GR_WR_DOUT[5]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i6.GSR = "DISABLED";
    CCU2D add_1840_3 (.A0(x[1]), .B0(x[2]), .C0(GND_net), .D0(GND_net), 
          .A1(x[2]), .B1(x[3]), .C1(GND_net), .D1(GND_net), .CIN(n14126), 
          .COUT(n14127), .S0(currAddress_17__N_742[2]), .S1(currAddress_17__N_742[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[150:167])
    defparam add_1840_3.INIT0 = 16'h5666;
    defparam add_1840_3.INIT1 = 16'h5666;
    defparam add_1840_3.INJECT1_0 = "NO";
    defparam add_1840_3.INJECT1_1 = "NO";
    PFUMX i13406 (.BLUT(n15403), .ALUT(n17264), .C0(state[7]), .Z(n17265));
    LUT4 i3_4_lut_4_lut_4_lut (.A(state[4]), .B(SpriteRead_xValid), .C(state[5]), 
         .D(\state[0] ), .Z(n14_adj_2075)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i3_4_lut_4_lut_4_lut.init = 16'h0008;
    MULT2 mult_9u_9u_0_mult_0_1_adj_359 (.A0(GREEN_READ[2]), .A1(GREEN_READ[3]), 
          .A2(GREEN_READ[3]), .A3(GREEN_READ[4]), .B0(ALPHA_READ[1]), 
          .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), 
          .CI(mco_adj_2078), .CO(mco_1_adj_2074), .P0(mult_9u_9u_0_pp_0_3_adj_2077), 
          .P1(mult_9u_9u_0_pp_0_4_adj_2076)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    MULT2 mult_9u_9u_0_mult_0_0_adj_360 (.A0(GREEN_READ[0]), .A1(GREEN_READ[1]), 
          .A2(GREEN_READ[1]), .A3(GREEN_READ[2]), .B0(ALPHA_READ[1]), 
          .B1(ALPHA_READ[0]), .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), 
          .CI(mult_9u_9u_0_cin_lr_0_adj_2011), .CO(mco_adj_2078), .P0(GREEN_OUT_9__N_669[1]), 
          .P1(mult_9u_9u_0_pp_0_2_adj_2079)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B t_mult_9u_9u_0_add_3_6_adj_361 (.A0(s_mult_9u_9u_0_2_17_adj_2081), 
           .A1(GND_net), .B0(GND_net), .B1(GND_net), .CI(co_t_mult_9u_9u_0_3_5_adj_2080), 
           .S0(GREEN_OUT_9__N_669[17])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 i22_3_lut_3_lut (.A(state[4]), .B(\state[0] ), .C(state[7]), 
         .Z(n11)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)+!B !(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i22_3_lut_3_lut.init = 16'h3434;
    LUT4 i13026_2_lut_rep_438 (.A(state[6]), .B(state[5]), .Z(n17446)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i13026_2_lut_rep_438.init = 16'h1111;
    LUT4 i12379_3_lut (.A(n3975), .B(n3991), .C(currSprite[4]), .Z(n16041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12379_3_lut.init = 16'hcaca;
    LUT4 i13068_2_lut_4_lut (.A(n1193), .B(n17361), .C(n17360), .D(n15_adj_2082), 
         .Z(LOGIC_CLOCK_enable_13)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (B+!(C (D))))) */ ;
    defparam i13068_2_lut_4_lut.init = 16'h3a00;
    LUT4 LED_c_bdd_2_lut_3_lut_13868 (.A(state[6]), .B(state[5]), .C(n17263), 
         .Z(n17264)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam LED_c_bdd_2_lut_3_lut_13868.init = 16'h1010;
    CCU2D BLUE_OUT_9__I_0_12 (.A0(BLUE_OUT_9__N_687[10]), .B0(BLUE_OUT_9__N_706[10]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[11]), .B1(BLUE_OUT_9__N_706[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14052), .COUT(n14053), .S0(BLUE_OUT[1]), 
          .S1(BLUE_OUT[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_12.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_12.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_12.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_12.INJECT1_1 = "NO";
    FADD2B t_mult_9u_9u_0_add_3_5_adj_362 (.A0(s_mult_9u_9u_0_2_15_adj_2084), 
           .A1(s_mult_9u_9u_0_2_16_adj_2085), .B0(mult_9u_9u_0_pp_4_15_adj_2013), 
           .B1(mult_9u_9u_0_pp_4_16_adj_2012), .CI(co_t_mult_9u_9u_0_3_4_adj_2083), 
           .COUT(co_t_mult_9u_9u_0_3_5_adj_2080), .S0(GREEN_OUT_9__N_669[15]), 
           .S1(GREEN_OUT_9__N_669[16])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B t_mult_9u_9u_0_add_3_4_adj_363 (.A0(s_mult_9u_9u_0_2_13_adj_2087), 
           .A1(s_mult_9u_9u_0_2_14_adj_2088), .B0(mult_9u_9u_0_pp_4_13_adj_2015), 
           .B1(mult_9u_9u_0_pp_4_14_adj_2014), .CI(co_t_mult_9u_9u_0_3_3_adj_2086), 
           .COUT(co_t_mult_9u_9u_0_3_4_adj_2083), .S0(GREEN_OUT_9__N_669[13]), 
           .S1(GREEN_OUT_9__N_669[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 n10147_bdd_4_lut_13400 (.A(n17396), .B(n17275), .C(n14447), .D(\state[1] ), 
         .Z(n17255)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam n10147_bdd_4_lut_13400.init = 16'h0511;
    FADD2B t_mult_9u_9u_0_add_3_3_adj_364 (.A0(s_mult_9u_9u_0_2_11_adj_2090), 
           .A1(s_mult_9u_9u_0_2_12_adj_2091), .B0(mult_9u_9u_0_pp_4_11_adj_2017), 
           .B1(mult_9u_9u_0_pp_4_12_adj_2016), .CI(co_t_mult_9u_9u_0_3_2_adj_2089), 
           .COUT(co_t_mult_9u_9u_0_3_3_adj_2086), .S0(GREEN_OUT_9__N_669[11]), 
           .S1(GREEN_OUT_9__N_669[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B t_mult_9u_9u_0_add_3_2_adj_365 (.A0(s_mult_9u_9u_0_2_9_adj_2093), 
           .A1(s_mult_9u_9u_0_2_10_adj_2094), .B0(mult_9u_9u_0_pp_4_9_adj_2019), 
           .B1(mult_9u_9u_0_pp_4_10_adj_2018), .CI(co_t_mult_9u_9u_0_3_1_adj_2092), 
           .COUT(co_t_mult_9u_9u_0_3_2_adj_2089), .S0(GREEN_OUT_9__N_669[9]), 
           .S1(GREEN_OUT_9__N_669[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B Cadd_t_mult_9u_9u_0_3_1_adj_366 (.A0(GND_net), .A1(s_mult_9u_9u_0_2_8_adj_2095), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_4_8_adj_1880), .CI(GND_net), 
           .COUT(co_t_mult_9u_9u_0_3_1_adj_2092), .S1(GREEN_OUT_9__N_669[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_2_8_adj_367 (.A0(GND_net), .A1(GND_net), .B0(s_mult_9u_9u_0_1_17_adj_2097), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_2_7_adj_2096), .S0(s_mult_9u_9u_0_2_17_adj_2081)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    CCU2D yPre_7__I_0_757_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(MATRIX_CURRROW[0]), .B1(yOffset[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n14016), .S1(currAddress_17__N_724[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[24:38])
    defparam yPre_7__I_0_757_1.INIT0 = 16'hF000;
    defparam yPre_7__I_0_757_1.INIT1 = 16'ha999;
    defparam yPre_7__I_0_757_1.INJECT1_0 = "NO";
    defparam yPre_7__I_0_757_1.INJECT1_1 = "NO";
    LUT4 i6587_2_lut_4_lut (.A(n23_adj_1904), .B(SpriteRead_xValid), .C(state[4]), 
         .D(\state[0] ), .Z(n9918)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i6587_2_lut_4_lut.init = 16'hffca;
    FADD2B mult_9u_9u_0_add_2_7_adj_368 (.A0(GND_net), .A1(GND_net), .B0(s_mult_9u_9u_0_1_15_adj_2099), 
           .B1(s_mult_9u_9u_0_1_16_adj_2100), .CI(co_mult_9u_9u_0_2_6_adj_2098), 
           .COUT(co_mult_9u_9u_0_2_7_adj_2096), .S0(s_mult_9u_9u_0_2_15_adj_2084), 
           .S1(s_mult_9u_9u_0_2_16_adj_2085)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_2_6_adj_369 (.A0(s_mult_9u_9u_0_0_13_adj_2104), 
           .A1(GND_net), .B0(s_mult_9u_9u_0_1_13_adj_2102), .B1(s_mult_9u_9u_0_1_14_adj_2103), 
           .CI(co_mult_9u_9u_0_2_5_adj_2101), .COUT(co_mult_9u_9u_0_2_6_adj_2098), 
           .S0(s_mult_9u_9u_0_2_13_adj_2087), .S1(s_mult_9u_9u_0_2_14_adj_2088)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_2_5_adj_370 (.A0(s_mult_9u_9u_0_0_11_adj_2108), 
           .A1(s_mult_9u_9u_0_0_12_adj_2109), .B0(s_mult_9u_9u_0_1_11_adj_2106), 
           .B1(s_mult_9u_9u_0_1_12_adj_2107), .CI(co_mult_9u_9u_0_2_4_adj_2105), 
           .COUT(co_mult_9u_9u_0_2_5_adj_2101), .S0(s_mult_9u_9u_0_2_11_adj_2090), 
           .S1(s_mult_9u_9u_0_2_12_adj_2091)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_2_4_adj_371 (.A0(s_mult_9u_9u_0_0_9_adj_2113), 
           .A1(s_mult_9u_9u_0_0_10_adj_2114), .B0(s_mult_9u_9u_0_1_9_adj_2111), 
           .B1(s_mult_9u_9u_0_1_10_adj_2112), .CI(co_mult_9u_9u_0_2_3_adj_2110), 
           .COUT(co_mult_9u_9u_0_2_4_adj_2105), .S0(s_mult_9u_9u_0_2_9_adj_2093), 
           .S1(s_mult_9u_9u_0_2_10_adj_2094)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_2_3_adj_372 (.A0(s_mult_9u_9u_0_0_7_adj_2118), 
           .A1(s_mult_9u_9u_0_0_8_adj_2119), .B0(s_mult_9u_9u_0_1_7_adj_2116), 
           .B1(s_mult_9u_9u_0_1_8_adj_2117), .CI(co_mult_9u_9u_0_2_2_adj_2115), 
           .COUT(co_mult_9u_9u_0_2_3_adj_2110), .S0(GREEN_OUT_9__N_669[7]), 
           .S1(s_mult_9u_9u_0_2_8_adj_2095)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_2_2 (.A0(s_mult_9u_9u_0_0_5_adj_2121), .A1(s_mult_9u_9u_0_0_6_adj_2122), 
           .B0(mult_9u_9u_0_pp_2_5_adj_2049), .B1(s_mult_9u_9u_0_1_6_adj_2120), 
           .CI(co_mult_9u_9u_0_2_1), .COUT(co_mult_9u_9u_0_2_2_adj_2115), 
           .S0(GREEN_OUT_9__N_669[5]), .S1(GREEN_OUT_9__N_669[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    PFUMX i12101 (.BLUT(n15761), .ALUT(n15762), .C0(n17334), .Z(Sprite_readData2_15__N_524[5]));
    LUT4 i2_3_lut_rep_388_4_lut (.A(state[6]), .B(state[5]), .C(state[4]), 
         .D(\state[3] ), .Z(n17396)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_388_4_lut.init = 16'hfffe;
    LUT4 i12989_2_lut_rep_398_3_lut (.A(state[6]), .B(state[5]), .C(\state[3] ), 
         .Z(n17406)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i12989_2_lut_rep_398_3_lut.init = 16'h0101;
    FADD2B Cadd_mult_9u_9u_0_2_1 (.A0(GND_net), .A1(s_mult_9u_9u_0_0_4_adj_2124), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_2_4_adj_2123), .CI(GND_net), 
           .COUT(co_mult_9u_9u_0_2_1), .S1(GREEN_OUT_9__N_669[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B Cadd_mult_9u_9u_0_1_7 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_1_6_adj_2125), .S0(s_mult_9u_9u_0_1_17_adj_2097)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_1_6_adj_373 (.A0(GND_net), .A1(GND_net), .B0(mult_9u_9u_0_pp_3_15_adj_2021), 
           .B1(mult_9u_9u_0_pp_3_16_adj_2020), .CI(co_mult_9u_9u_0_1_5_adj_2126), 
           .COUT(co_mult_9u_9u_0_1_6_adj_2125), .S0(s_mult_9u_9u_0_1_15_adj_2099), 
           .S1(s_mult_9u_9u_0_1_16_adj_2100)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_1_5_adj_374 (.A0(mult_9u_9u_0_pp_2_13_adj_2037), 
           .A1(mult_9u_9u_0_pp_2_14_adj_2036), .B0(mult_9u_9u_0_pp_3_13_adj_2025), 
           .B1(mult_9u_9u_0_pp_3_14_adj_2024), .CI(co_mult_9u_9u_0_1_4_adj_2127), 
           .COUT(co_mult_9u_9u_0_1_5_adj_2126), .S0(s_mult_9u_9u_0_1_13_adj_2102), 
           .S1(s_mult_9u_9u_0_1_14_adj_2103)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_1_4_adj_375 (.A0(mult_9u_9u_0_pp_2_11_adj_2040), 
           .A1(mult_9u_9u_0_pp_2_12_adj_2039), .B0(mult_9u_9u_0_pp_3_11_adj_2028), 
           .B1(mult_9u_9u_0_pp_3_12_adj_2027), .CI(co_mult_9u_9u_0_1_3_adj_2128), 
           .COUT(co_mult_9u_9u_0_1_4_adj_2127), .S0(s_mult_9u_9u_0_1_11_adj_2106), 
           .S1(s_mult_9u_9u_0_1_12_adj_2107)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 i257_2_lut_rep_263_2_lut (.A(n17275), .B(n1), .Z(n17271)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i257_2_lut_rep_263_2_lut.init = 16'h1111;
    LUT4 i1_2_lut (.A(state[7]), .B(state[6]), .Z(n15442)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i12991_3_lut (.A(n15701), .B(MATRIX_CURRROW[0]), .C(n15_adj_2023), 
         .Z(LOGIC_CLOCK_enable_50)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam i12991_3_lut.init = 16'h0202;
    FADD2B mult_9u_9u_0_add_1_3_adj_376 (.A0(mult_9u_9u_0_pp_2_9_adj_2043), 
           .A1(mult_9u_9u_0_pp_2_10_adj_2042), .B0(mult_9u_9u_0_pp_3_9_adj_2031), 
           .B1(mult_9u_9u_0_pp_3_10_adj_2030), .CI(co_mult_9u_9u_0_1_2_adj_2129), 
           .COUT(co_mult_9u_9u_0_1_3_adj_2128), .S0(s_mult_9u_9u_0_1_9_adj_2111), 
           .S1(s_mult_9u_9u_0_1_10_adj_2112)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_1_2_adj_377 (.A0(mult_9u_9u_0_pp_2_7_adj_2046), 
           .A1(mult_9u_9u_0_pp_2_8_adj_2045), .B0(mult_9u_9u_0_pp_3_7_adj_2034), 
           .B1(mult_9u_9u_0_pp_3_8_adj_2033), .CI(co_mult_9u_9u_0_1_1_adj_2130), 
           .COUT(co_mult_9u_9u_0_1_2_adj_2129), .S0(s_mult_9u_9u_0_1_7_adj_2116), 
           .S1(s_mult_9u_9u_0_1_8_adj_2117)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B Cadd_mult_9u_9u_0_1_1_adj_378 (.A0(GND_net), .A1(mult_9u_9u_0_pp_2_6_adj_2048), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_3_6_adj_2131), .CI(GND_net), 
           .COUT(co_mult_9u_9u_0_1_1_adj_2130), .S1(s_mult_9u_9u_0_1_6_adj_2120)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B Cadd_mult_9u_9u_0_0_7_adj_379 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_0_6_adj_2132), .S0(s_mult_9u_9u_0_0_13_adj_2104)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_0_6_adj_380 (.A0(GND_net), .A1(GND_net), .B0(mult_9u_9u_0_pp_1_11_adj_2052), 
           .B1(mult_9u_9u_0_pp_1_12_adj_2051), .CI(co_mult_9u_9u_0_0_5_adj_2133), 
           .COUT(co_mult_9u_9u_0_0_6_adj_2132), .S0(s_mult_9u_9u_0_0_11_adj_2108), 
           .S1(s_mult_9u_9u_0_0_12_adj_2109)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_0_5_adj_381 (.A0(mult_9u_9u_0_pp_0_9_adj_2067), 
           .A1(mult_9u_9u_0_pp_0_10_adj_2066), .B0(mult_9u_9u_0_pp_1_9_adj_2055), 
           .B1(mult_9u_9u_0_pp_1_10_adj_2054), .CI(co_mult_9u_9u_0_0_4_adj_2134), 
           .COUT(co_mult_9u_9u_0_0_5_adj_2133), .S0(s_mult_9u_9u_0_0_9_adj_2113), 
           .S1(s_mult_9u_9u_0_0_10_adj_2114)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_0_4_adj_382 (.A0(mult_9u_9u_0_pp_0_7_adj_2070), 
           .A1(mult_9u_9u_0_pp_0_8_adj_2069), .B0(mult_9u_9u_0_pp_1_7_adj_2058), 
           .B1(mult_9u_9u_0_pp_1_8_adj_2057), .CI(co_mult_9u_9u_0_0_3_adj_2135), 
           .COUT(co_mult_9u_9u_0_0_4_adj_2134), .S0(s_mult_9u_9u_0_0_7_adj_2118), 
           .S1(s_mult_9u_9u_0_0_8_adj_2119)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    LUT4 i12040_4_lut (.A(MATRIX_CURRROW[2]), .B(MATRIX_CURRROW[1]), .C(MATRIX_CURRROW[3]), 
         .D(MATRIX_CURRROW[4]), .Z(n15701)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12040_4_lut.init = 16'h8000;
    FD1P3AX GR_WR_DOUT_16__i5 (.D(GR_WR_DOUT[4]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i5.GSR = "DISABLED";
    FD1P3AX GR_WR_DOUT_16__i4 (.D(GR_WR_DOUT[3]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i4.GSR = "DISABLED";
    FD1P3AX GR_WR_DOUT_16__i3 (.D(GR_WR_DOUT[2]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i3.GSR = "DISABLED";
    LUT4 i12378_3_lut (.A(n3940), .B(n3956), .C(currSprite[4]), .Z(n16040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12378_3_lut.init = 16'hcaca;
    FADD2B mult_9u_9u_0_add_0_3_adj_383 (.A0(mult_9u_9u_0_pp_0_5_adj_2073), 
           .A1(mult_9u_9u_0_pp_0_6_adj_2072), .B0(mult_9u_9u_0_pp_1_5_adj_2061), 
           .B1(mult_9u_9u_0_pp_1_6_adj_2060), .CI(co_mult_9u_9u_0_0_2_adj_2136), 
           .COUT(co_mult_9u_9u_0_0_3_adj_2135), .S0(s_mult_9u_9u_0_0_5_adj_2121), 
           .S1(s_mult_9u_9u_0_0_6_adj_2122)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_add_0_2_adj_384 (.A0(mult_9u_9u_0_pp_0_3_adj_2077), 
           .A1(mult_9u_9u_0_pp_0_4_adj_2076), .B0(mult_9u_9u_0_pp_1_3_adj_2064), 
           .B1(mult_9u_9u_0_pp_1_4_adj_2063), .CI(co_mult_9u_9u_0_0_1_adj_2137), 
           .COUT(co_mult_9u_9u_0_0_2_adj_2136), .S0(GREEN_OUT_9__N_669[3]), 
           .S1(s_mult_9u_9u_0_0_4_adj_2124)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B Cadd_mult_9u_9u_0_0_1_adj_385 (.A0(GND_net), .A1(mult_9u_9u_0_pp_0_2_adj_2079), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_1_2_adj_2138), .CI(GND_net), 
           .COUT(co_mult_9u_9u_0_0_1_adj_2137), .S1(GREEN_OUT_9__N_669[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_cin_lr_add_6_adj_386 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_6_adj_2035)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_cin_lr_add_4_adj_387 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_4_adj_2050)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FADD2B mult_9u_9u_0_cin_lr_add_2_adj_388 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_2_adj_2065)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[132:152])
    FD1P3AX GR_WR_DOUT_16__i2 (.D(GR_WR_DOUT[1]), .SP(LOGIC_CLOCK_enable_79), 
            .CK(LOGIC_CLOCK), .Q(GR_WR_DOUT_16[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam GR_WR_DOUT_16__i2.GSR = "DISABLED";
    PFUMX i12562 (.BLUT(n16216), .ALUT(n16217), .C0(n17334), .Z(n16224));
    LUT4 i1_2_lut_rep_361_3_lut_4_lut (.A(state[6]), .B(state[5]), .C(\state[1] ), 
         .D(\state[3] ), .Z(n17369)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_361_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12376_3_lut (.A(n3973), .B(n3989), .C(currSprite[4]), .Z(n16038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12376_3_lut.init = 16'hcaca;
    CCU2D xPre_7__I_0_752_8 (.A0(xPre[6]), .B0(xOffset_c[6]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[7]), .B1(xOffset_c[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14014), .S0(x[6]), .S1(x[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(249[25:39])
    defparam xPre_7__I_0_752_8.INIT0 = 16'h5666;
    defparam xPre_7__I_0_752_8.INIT1 = 16'h5666;
    defparam xPre_7__I_0_752_8.INJECT1_0 = "NO";
    defparam xPre_7__I_0_752_8.INJECT1_1 = "NO";
    AND2 AND2_t12_adj_389 (.A(GREEN_READ[0]), .B(ALPHA_READ[0]), .Z(GREEN_OUT_9__N_669[0])) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(159[10:64])
    LUT4 i12375_3_lut (.A(n3938), .B(n3954), .C(currSprite[4]), .Z(n16037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12375_3_lut.init = 16'hcaca;
    PFUMX i12563 (.BLUT(n16218), .ALUT(n16219), .C0(n17334), .Z(n16225));
    AND2 AND2_t11_adj_390 (.A(GREEN_READ[0]), .B(ALPHA_READ[2]), .Z(mult_9u_9u_0_pp_1_2_adj_2138)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(161[10:64])
    LUT4 i12373_3_lut (.A(n3962), .B(n3978), .C(currSprite[4]), .Z(n16035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12373_3_lut.init = 16'hcaca;
    LUT4 i928_3_lut_4_lut (.A(state[4]), .B(SpriteRead_xValid), .C(n8625), 
         .D(\state[0] ), .Z(n3201)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i928_3_lut_4_lut.init = 16'h8f88;
    PFUMX i12564 (.BLUT(n16220), .ALUT(n16221), .C0(n17334), .Z(n16226));
    FADD2B mult_9u_9u_0_add_2_2_adj_391 (.A0(s_mult_9u_9u_0_0_5), .A1(s_mult_9u_9u_0_0_6), 
           .B0(mult_9u_9u_0_pp_2_5), .B1(s_mult_9u_9u_0_1_6), .CI(co_mult_9u_9u_0_2_1_adj_2139), 
           .COUT(co_mult_9u_9u_0_2_2), .S0(RED_OUT_9__N_632[5]), .S1(RED_OUT_9__N_632[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    AND2 AND2_t10_adj_392 (.A(GREEN_READ[0]), .B(ALPHA_READ[4]), .Z(mult_9u_9u_0_pp_2_4_adj_2123)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(163[10:64])
    AND2 AND2_t9_adj_393 (.A(GREEN_READ[0]), .B(ALPHA_READ[6]), .Z(mult_9u_9u_0_pp_3_6_adj_2131)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(165[10:63])
    FADD2B mult_10u_9u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    AND2 AND2_t0_adj_394 (.A(VRAM_DATA_OUT[19]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_17)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(196[10:65])
    AND2 AND2_t1_adj_395 (.A(VRAM_DATA_OUT[18]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(194[10:65])
    AND2 AND2_t2_adj_396 (.A(VRAM_DATA_OUT[17]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_15)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(192[10:65])
    AND2 AND2_t9_adj_397 (.A(VRAM_DATA_OUT[0]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_8_adj_2140)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(178[10:64])
    LUT4 i12372_3_lut (.A(n3927), .B(n3943), .C(currSprite[4]), .Z(n16034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12372_3_lut.init = 16'hcaca;
    AND2 AND2_t3_adj_398 (.A(VRAM_DATA_OUT[16]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(190[10:65])
    AND2 AND2_t4_adj_399 (.A(VRAM_DATA_OUT[15]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_13)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(188[10:65])
    AND2 AND2_t5_adj_400 (.A(VRAM_DATA_OUT[14]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(186[10:65])
    AND2 AND2_t6_adj_401 (.A(VRAM_DATA_OUT[13]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_11)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(184[10:65])
    AND2 AND2_t7_adj_402 (.A(VRAM_DATA_OUT[12]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(182[10:65])
    AND2 AND2_t8_adj_403 (.A(VRAM_DATA_OUT[11]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_9)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(180[10:64])
    PFUMX i13404 (.BLUT(n17262), .ALUT(n15343), .C0(state[4]), .Z(n17263));
    PFUMX i12565 (.BLUT(n16222), .ALUT(n16223), .C0(n17334), .Z(n16227));
    LUT4 i1_2_lut_3_lut_4_lut_adj_404 (.A(state[6]), .B(state[5]), .C(state[4]), 
         .D(\state[3] ), .Z(n4_adj_2141)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_404.init = 16'h0010;
    MULT2 mult_10u_9u_0_mult_6_4 (.A0(VRAM_DATA_OUT[18]), .A1(VRAM_DATA_OUT[19]), 
          .A2(VRAM_DATA_OUT[19]), .A3(GND_net), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_15_adj_2142), .CO(mfco_3), .P0(mult_10u_9u_0_pp_3_15), 
          .P1(mult_10u_9u_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_6_3 (.A0(VRAM_DATA_OUT[16]), .A1(VRAM_DATA_OUT[17]), 
          .A2(VRAM_DATA_OUT[17]), .A3(VRAM_DATA_OUT[18]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_14_adj_2143), .CO(mco_15_adj_2142), .P0(mult_10u_9u_0_pp_3_13), 
          .P1(mult_10u_9u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_6_2 (.A0(VRAM_DATA_OUT[14]), .A1(VRAM_DATA_OUT[15]), 
          .A2(VRAM_DATA_OUT[15]), .A3(VRAM_DATA_OUT[16]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_13_adj_2144), .CO(mco_14_adj_2143), .P0(mult_10u_9u_0_pp_3_11), 
          .P1(mult_10u_9u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_6_1 (.A0(VRAM_DATA_OUT[12]), .A1(VRAM_DATA_OUT[13]), 
          .A2(VRAM_DATA_OUT[13]), .A3(VRAM_DATA_OUT[14]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_12_adj_2145), .CO(mco_13_adj_2144), .P0(mult_10u_9u_0_pp_3_9), 
          .P1(mult_10u_9u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_6_0 (.A0(VRAM_DATA_OUT[10]), .A1(VRAM_DATA_OUT[11]), 
          .A2(VRAM_DATA_OUT[11]), .A3(VRAM_DATA_OUT[12]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mult_10u_9u_0_cin_lr_6), .CO(mco_12_adj_2145), .P0(mult_10u_9u_0_pp_3_7), 
          .P1(mult_10u_9u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    FD1P3AX reset_706 (.D(reset_N_1062), .SP(state_7__N_345), .CK(LOGIC_CLOCK), 
            .Q(reset)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam reset_706.GSR = "DISABLED";
    FADD2B Cadd_mult_9u_9u_0_2_1_adj_405 (.A0(GND_net), .A1(s_mult_9u_9u_0_0_4), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_2_4), .CI(GND_net), .COUT(co_mult_9u_9u_0_2_1_adj_2139), 
           .S1(RED_OUT_9__N_632[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    MULT2 mult_10u_9u_0_mult_4_4 (.A0(VRAM_DATA_OUT[18]), .A1(VRAM_DATA_OUT[19]), 
          .A2(VRAM_DATA_OUT[19]), .A3(GND_net), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_11_adj_2146), .CO(mfco_2), .P0(mult_10u_9u_0_pp_2_13), 
          .P1(mult_10u_9u_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_4_3 (.A0(VRAM_DATA_OUT[16]), .A1(VRAM_DATA_OUT[17]), 
          .A2(VRAM_DATA_OUT[17]), .A3(VRAM_DATA_OUT[18]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_10_adj_2147), .CO(mco_11_adj_2146), .P0(mult_10u_9u_0_pp_2_11), 
          .P1(mult_10u_9u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_4_2 (.A0(VRAM_DATA_OUT[14]), .A1(VRAM_DATA_OUT[15]), 
          .A2(VRAM_DATA_OUT[15]), .A3(VRAM_DATA_OUT[16]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_9_adj_2148), .CO(mco_10_adj_2147), .P0(mult_10u_9u_0_pp_2_9), 
          .P1(mult_10u_9u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_4_1 (.A0(VRAM_DATA_OUT[12]), .A1(VRAM_DATA_OUT[13]), 
          .A2(VRAM_DATA_OUT[13]), .A3(VRAM_DATA_OUT[14]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_8_adj_2149), .CO(mco_9_adj_2148), .P0(mult_10u_9u_0_pp_2_7), 
          .P1(mult_10u_9u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_4_0 (.A0(VRAM_DATA_OUT[10]), .A1(VRAM_DATA_OUT[11]), 
          .A2(VRAM_DATA_OUT[11]), .A3(VRAM_DATA_OUT[12]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mult_10u_9u_0_cin_lr_4), .CO(mco_8_adj_2149), .P0(mult_10u_9u_0_pp_2_5), 
          .P1(mult_10u_9u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    CCU2D add_1840_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[0]), .B1(xOffset[0]), .C1(x[1]), .D1(GND_net), .COUT(n14126), 
          .S1(currAddress_17__N_742[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[150:167])
    defparam add_1840_1.INIT0 = 16'hF000;
    defparam add_1840_1.INIT1 = 16'h9696;
    defparam add_1840_1.INJECT1_0 = "NO";
    defparam add_1840_1.INJECT1_1 = "NO";
    FD1P3AX Sprite_writeClk_740 (.D(Sprite_writeClk_N_1144), .SP(LOGIC_CLOCK_enable_81), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeClk)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeClk_740.GSR = "DISABLED";
    CCU2D add_10518_15 (.A0(n16[13]), .B0(\Sprite_readAddr_13__N_752[13] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14125), .S0(Sprite_readAddr[13]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_15.INIT0 = 16'h5666;
    defparam add_10518_15.INIT1 = 16'h0000;
    defparam add_10518_15.INJECT1_0 = "NO";
    defparam add_10518_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_406 (.A(n17458), .B(n17329), .C(n17313), 
         .D(n17273), .Z(n3960)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(570[10:40])
    defparam i1_2_lut_3_lut_4_lut_adj_406.init = 16'h0200;
    LUT4 i12370_3_lut (.A(n3970), .B(n3986), .C(currSprite[4]), .Z(n16032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12370_3_lut.init = 16'hcaca;
    CCU2D add_10518_13 (.A0(n16[11]), .B0(\Sprite_readAddr_13__N_752[11] ), 
          .C0(GND_net), .D0(GND_net), .A1(n16[12]), .B1(\Sprite_readAddr_13__N_752[12] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14124), .COUT(n14125), .S0(Sprite_readAddr[11]), 
          .S1(Sprite_readAddr[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_13.INIT0 = 16'h5666;
    defparam add_10518_13.INIT1 = 16'h5666;
    defparam add_10518_13.INJECT1_0 = "NO";
    defparam add_10518_13.INJECT1_1 = "NO";
    CCU2D add_10518_11 (.A0(n16[9]), .B0(\Sprite_readAddr_13__N_752[9] ), 
          .C0(GND_net), .D0(GND_net), .A1(n16[10]), .B1(\Sprite_readAddr_13__N_752[10] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14123), .COUT(n14124), .S0(Sprite_readAddr[9]), 
          .S1(Sprite_readAddr[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_11.INIT0 = 16'h5666;
    defparam add_10518_11.INIT1 = 16'h5666;
    defparam add_10518_11.INJECT1_0 = "NO";
    defparam add_10518_11.INJECT1_1 = "NO";
    MULT2 mult_10u_9u_0_mult_2_4 (.A0(VRAM_DATA_OUT[18]), .A1(VRAM_DATA_OUT[19]), 
          .A2(VRAM_DATA_OUT[19]), .A3(GND_net), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_7_adj_2150), .CO(mfco_1), .P0(mult_10u_9u_0_pp_1_11), 
          .P1(mult_10u_9u_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    LUT4 i1_4_lut_4_lut_adj_407 (.A(SpriteRead_xValid), .B(n70), .C(state[2]), 
         .D(n15699), .Z(n15343)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_adj_407.init = 16'h00f4;
    PFUMX i13416 (.BLUT(n17483), .ALUT(n17484), .C0(state[4]), .Z(n17485));
    LUT4 i6907_3_lut_4_lut_4_lut (.A(n17275), .B(SpriteRead_yInSprite_7__N_597[5]), 
         .C(n17318), .D(n1), .Z(n2191[0])) /* synthesis lut_function=(A (B (C))+!A (B (C (D))+!B !((D)+!C))) */ ;
    defparam i6907_3_lut_4_lut_4_lut.init = 16'hc090;
    LUT4 i2_4_lut_adj_408 (.A(n17276), .B(BUS_transferState[2]), .C(n17), 
         .D(LOGIC_CLOCK_enable_52), .Z(n15352)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[4] 608[11])
    defparam i2_4_lut_adj_408.init = 16'h0010;
    MULT2 mult_10u_9u_0_mult_2_3 (.A0(VRAM_DATA_OUT[16]), .A1(VRAM_DATA_OUT[17]), 
          .A2(VRAM_DATA_OUT[17]), .A3(VRAM_DATA_OUT[18]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_6_adj_2151), .CO(mco_7_adj_2150), .P0(mult_10u_9u_0_pp_1_9), 
          .P1(mult_10u_9u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_2_2 (.A0(VRAM_DATA_OUT[14]), .A1(VRAM_DATA_OUT[15]), 
          .A2(VRAM_DATA_OUT[15]), .A3(VRAM_DATA_OUT[16]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_5_adj_2152), .CO(mco_6_adj_2151), .P0(mult_10u_9u_0_pp_1_7), 
          .P1(mult_10u_9u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_2_1 (.A0(VRAM_DATA_OUT[12]), .A1(VRAM_DATA_OUT[13]), 
          .A2(VRAM_DATA_OUT[13]), .A3(VRAM_DATA_OUT[14]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_4_adj_2153), .CO(mco_5_adj_2152), .P0(mult_10u_9u_0_pp_1_5), 
          .P1(mult_10u_9u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    MULT2 mult_10u_9u_0_mult_2_0 (.A0(VRAM_DATA_OUT[10]), .A1(VRAM_DATA_OUT[11]), 
          .A2(VRAM_DATA_OUT[11]), .A3(VRAM_DATA_OUT[12]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mult_10u_9u_0_cin_lr_2), .CO(mco_4_adj_2153), .P0(mult_10u_9u_0_pp_1_3), 
          .P1(mult_10u_9u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[61:103])
    PFUMX i12104 (.BLUT(n15764), .ALUT(n15765), .C0(n17334), .Z(Sprite_readData2_15__N_524[6]));
    LUT4 i12369_3_lut (.A(n3935), .B(n3951), .C(currSprite[4]), .Z(n16031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12369_3_lut.init = 16'hcaca;
    FADD2B Cadd_mult_9u_9u_0_1_7_adj_409 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_1_6), .S0(s_mult_9u_9u_0_1_17)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[126:146])
    FADD2B mult_10u_9u_0_add_2_5_adj_410 (.A0(s_mult_10u_9u_0_0_11_adj_1968), 
           .A1(s_mult_10u_9u_0_0_12_adj_1969), .B0(s_mult_10u_9u_0_1_11_adj_1940), 
           .B1(s_mult_10u_9u_0_1_12_adj_1941), .CI(co_mult_10u_9u_0_2_4_adj_2154), 
           .COUT(co_mult_10u_9u_0_2_5_adj_1909), .S0(s_mult_10u_9u_0_2_11_adj_2155), 
           .S1(s_mult_10u_9u_0_2_12_adj_2156)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_2_4_adj_411 (.A0(s_mult_10u_9u_0_0_9_adj_1973), 
           .A1(s_mult_10u_9u_0_0_10_adj_1974), .B0(s_mult_10u_9u_0_1_9_adj_1947), 
           .B1(s_mult_10u_9u_0_1_10_adj_1948), .CI(co_mult_10u_9u_0_2_3_adj_2157), 
           .COUT(co_mult_10u_9u_0_2_4_adj_2154), .S0(s_mult_10u_9u_0_2_9_adj_2158), 
           .S1(s_mult_10u_9u_0_2_10_adj_2159)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_2_3_adj_412 (.A0(s_mult_10u_9u_0_0_7_adj_1980), 
           .A1(s_mult_10u_9u_0_0_8_adj_1981), .B0(s_mult_10u_9u_0_1_7_adj_1954), 
           .B1(s_mult_10u_9u_0_1_8_adj_1955), .CI(co_mult_10u_9u_0_2_2_adj_2160), 
           .COUT(co_mult_10u_9u_0_2_3_adj_2157), .S0(BLUE_OUT_9__N_687[7]), 
           .S1(s_mult_10u_9u_0_2_8_adj_2161)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B mult_10u_9u_0_add_2_2_adj_413 (.A0(s_mult_10u_9u_0_0_5_adj_1987), 
           .A1(s_mult_10u_9u_0_0_6_adj_1988), .B0(mult_10u_9u_0_pp_2_5_adj_2163), 
           .B1(s_mult_10u_9u_0_1_6_adj_1961), .CI(co_mult_10u_9u_0_2_1_adj_2162), 
           .COUT(co_mult_10u_9u_0_2_2_adj_2160), .S0(BLUE_OUT_9__N_687[5]), 
           .S1(BLUE_OUT_9__N_687[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B Cadd_mult_10u_9u_0_2_1_adj_414 (.A0(GND_net), .A1(s_mult_10u_9u_0_0_4_adj_1994), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_2_4_adj_2010), .CI(GND_net), 
           .COUT(co_mult_10u_9u_0_2_1_adj_2162), .S1(BLUE_OUT_9__N_687[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B Cadd_t_mult_10u_9u_0_3_1_adj_415 (.A0(GND_net), .A1(s_mult_10u_9u_0_2_8_adj_2161), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_4_8_adj_1881), .CI(GND_net), 
           .COUT(co_t_mult_10u_9u_0_3_1_adj_2164), .S1(BLUE_OUT_9__N_687[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B t_mult_10u_9u_0_add_3_2_adj_416 (.A0(s_mult_10u_9u_0_2_9_adj_2158), 
           .A1(s_mult_10u_9u_0_2_10_adj_2159), .B0(mult_10u_9u_0_pp_4_9_adj_2165), 
           .B1(mult_10u_9u_0_pp_4_10_adj_2166), .CI(co_t_mult_10u_9u_0_3_1_adj_2164), 
           .COUT(co_t_mult_10u_9u_0_3_2_adj_2167), .S0(BLUE_OUT_9__N_687[9]), 
           .S1(BLUE_OUT_9__N_687[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B t_mult_10u_9u_0_add_3_3_adj_417 (.A0(s_mult_10u_9u_0_2_11_adj_2155), 
           .A1(s_mult_10u_9u_0_2_12_adj_2156), .B0(mult_10u_9u_0_pp_4_11_adj_2168), 
           .B1(mult_10u_9u_0_pp_4_12_adj_2169), .CI(co_t_mult_10u_9u_0_3_2_adj_2167), 
           .COUT(co_t_mult_10u_9u_0_3_3_adj_2170), .S0(BLUE_OUT_9__N_687[11]), 
           .S1(BLUE_OUT_9__N_687[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B t_mult_10u_9u_0_add_3_4_adj_418 (.A0(s_mult_10u_9u_0_2_13_adj_1915), 
           .A1(s_mult_10u_9u_0_2_14_adj_1916), .B0(mult_10u_9u_0_pp_4_13_adj_2171), 
           .B1(mult_10u_9u_0_pp_4_14_adj_2172), .CI(co_t_mult_10u_9u_0_3_3_adj_2170), 
           .COUT(co_t_mult_10u_9u_0_3_4_adj_2173), .S0(BLUE_OUT_9__N_687[13]), 
           .S1(BLUE_OUT_9__N_687[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B t_mult_10u_9u_0_add_3_5_adj_419 (.A0(s_mult_10u_9u_0_2_15_adj_1922), 
           .A1(s_mult_10u_9u_0_2_16_adj_1923), .B0(mult_10u_9u_0_pp_4_15_adj_2174), 
           .B1(mult_10u_9u_0_pp_4_16_adj_2175), .CI(co_t_mult_10u_9u_0_3_4_adj_2173), 
           .COUT(co_t_mult_10u_9u_0_3_5_adj_2176), .S0(BLUE_OUT_9__N_687[15]), 
           .S1(BLUE_OUT_9__N_687[16])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    FADD2B t_mult_10u_9u_0_add_3_6_adj_420 (.A0(s_mult_10u_9u_0_2_17_adj_1926), 
           .A1(s_mult_10u_9u_0_2_18_adj_1927), .B0(mult_10u_9u_0_pp_4_17_adj_2177), 
           .B1(GND_net), .CI(co_t_mult_10u_9u_0_3_5_adj_2176), .S0(BLUE_OUT_9__N_687[17]), 
           .S1(BLUE_OUT_9__N_687[18])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_0_0_adj_421 (.A0(VRAM_DATA_OUT[20]), .A1(VRAM_DATA_OUT[21]), 
          .A2(VRAM_DATA_OUT[21]), .A3(VRAM_DATA_OUT[22]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mult_10u_9u_0_cin_lr_0_adj_2178), .CO(mco_adj_2179), .P0(BLUE_OUT_9__N_687[1]), 
          .P1(mult_10u_9u_0_pp_0_2_adj_2000)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_0_1_adj_422 (.A0(VRAM_DATA_OUT[22]), .A1(VRAM_DATA_OUT[23]), 
          .A2(VRAM_DATA_OUT[23]), .A3(VRAM_DATA_OUT[24]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_adj_2179), .CO(mco_1_adj_2180), .P0(mult_10u_9u_0_pp_0_3_adj_1996), 
          .P1(mult_10u_9u_0_pp_0_4_adj_1995)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_0_2_adj_423 (.A0(VRAM_DATA_OUT[24]), .A1(VRAM_DATA_OUT[25]), 
          .A2(VRAM_DATA_OUT[25]), .A3(VRAM_DATA_OUT[26]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_1_adj_2180), .CO(mco_2_adj_2181), .P0(mult_10u_9u_0_pp_0_5_adj_1990), 
          .P1(mult_10u_9u_0_pp_0_6_adj_1989)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_0_3_adj_424 (.A0(VRAM_DATA_OUT[26]), .A1(VRAM_DATA_OUT[27]), 
          .A2(VRAM_DATA_OUT[27]), .A3(VRAM_DATA_OUT[28]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_2_adj_2181), .CO(mco_3_adj_2182), .P0(mult_10u_9u_0_pp_0_7_adj_1983), 
          .P1(mult_10u_9u_0_pp_0_8_adj_1982)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_0_4_adj_425 (.A0(VRAM_DATA_OUT[28]), .A1(VRAM_DATA_OUT[29]), 
          .A2(VRAM_DATA_OUT[29]), .A3(GND_net), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_3_adj_2182), .CO(mfco_adj_2009), .P0(mult_10u_9u_0_pp_0_9_adj_1976), 
          .P1(mult_10u_9u_0_pp_0_10_adj_1975)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_2_0_adj_426 (.A0(VRAM_DATA_OUT[20]), .A1(VRAM_DATA_OUT[21]), 
          .A2(VRAM_DATA_OUT[21]), .A3(VRAM_DATA_OUT[22]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mult_10u_9u_0_cin_lr_2_adj_2008), .CO(mco_4_adj_2183), .P0(mult_10u_9u_0_pp_1_3_adj_1998), 
          .P1(mult_10u_9u_0_pp_1_4_adj_1997)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_2_1_adj_427 (.A0(VRAM_DATA_OUT[22]), .A1(VRAM_DATA_OUT[23]), 
          .A2(VRAM_DATA_OUT[23]), .A3(VRAM_DATA_OUT[24]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_4_adj_2183), .CO(mco_5_adj_2184), .P0(mult_10u_9u_0_pp_1_5_adj_1992), 
          .P1(mult_10u_9u_0_pp_1_6_adj_1991)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_2_2_adj_428 (.A0(VRAM_DATA_OUT[24]), .A1(VRAM_DATA_OUT[25]), 
          .A2(VRAM_DATA_OUT[25]), .A3(VRAM_DATA_OUT[26]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_5_adj_2184), .CO(mco_6_adj_2185), .P0(mult_10u_9u_0_pp_1_7_adj_1985), 
          .P1(mult_10u_9u_0_pp_1_8_adj_1984)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_2_3_adj_429 (.A0(VRAM_DATA_OUT[26]), .A1(VRAM_DATA_OUT[27]), 
          .A2(VRAM_DATA_OUT[27]), .A3(VRAM_DATA_OUT[28]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_6_adj_2185), .CO(mco_7_adj_2186), .P0(mult_10u_9u_0_pp_1_9_adj_1978), 
          .P1(mult_10u_9u_0_pp_1_10_adj_1977)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_2_4_adj_430 (.A0(VRAM_DATA_OUT[28]), .A1(VRAM_DATA_OUT[29]), 
          .A2(VRAM_DATA_OUT[29]), .A3(GND_net), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_7_adj_2186), .CO(mfco_1_adj_2007), .P0(mult_10u_9u_0_pp_1_11_adj_1971), 
          .P1(mult_10u_9u_0_pp_1_12_adj_1970)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_4_0_adj_431 (.A0(VRAM_DATA_OUT[20]), .A1(VRAM_DATA_OUT[21]), 
          .A2(VRAM_DATA_OUT[21]), .A3(VRAM_DATA_OUT[22]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mult_10u_9u_0_cin_lr_4_adj_2006), .CO(mco_8_adj_2187), .P0(mult_10u_9u_0_pp_2_5_adj_2163), 
          .P1(mult_10u_9u_0_pp_2_6_adj_1962)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_4_1_adj_432 (.A0(VRAM_DATA_OUT[22]), .A1(VRAM_DATA_OUT[23]), 
          .A2(VRAM_DATA_OUT[23]), .A3(VRAM_DATA_OUT[24]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_8_adj_2187), .CO(mco_9_adj_2188), .P0(mult_10u_9u_0_pp_2_7_adj_1957), 
          .P1(mult_10u_9u_0_pp_2_8_adj_1956)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_4_2_adj_433 (.A0(VRAM_DATA_OUT[24]), .A1(VRAM_DATA_OUT[25]), 
          .A2(VRAM_DATA_OUT[25]), .A3(VRAM_DATA_OUT[26]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_9_adj_2188), .CO(mco_10_adj_2189), .P0(mult_10u_9u_0_pp_2_9_adj_1950), 
          .P1(mult_10u_9u_0_pp_2_10_adj_1949)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_4_3_adj_434 (.A0(VRAM_DATA_OUT[26]), .A1(VRAM_DATA_OUT[27]), 
          .A2(VRAM_DATA_OUT[27]), .A3(VRAM_DATA_OUT[28]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_10_adj_2189), .CO(mco_11_adj_2190), .P0(mult_10u_9u_0_pp_2_11_adj_1943), 
          .P1(mult_10u_9u_0_pp_2_12_adj_1942)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_4_4_adj_435 (.A0(VRAM_DATA_OUT[28]), .A1(VRAM_DATA_OUT[29]), 
          .A2(VRAM_DATA_OUT[29]), .A3(GND_net), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_11_adj_2190), .CO(mfco_2_adj_2003), .P0(mult_10u_9u_0_pp_2_13_adj_1936), 
          .P1(mult_10u_9u_0_pp_2_14_adj_1935)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_6_0_adj_436 (.A0(VRAM_DATA_OUT[20]), .A1(VRAM_DATA_OUT[21]), 
          .A2(VRAM_DATA_OUT[21]), .A3(VRAM_DATA_OUT[22]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mult_10u_9u_0_cin_lr_6_adj_2002), .CO(mco_12_adj_2191), .P0(mult_10u_9u_0_pp_3_7_adj_1959), 
          .P1(mult_10u_9u_0_pp_3_8_adj_1958)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_6_1_adj_437 (.A0(VRAM_DATA_OUT[22]), .A1(VRAM_DATA_OUT[23]), 
          .A2(VRAM_DATA_OUT[23]), .A3(VRAM_DATA_OUT[24]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_12_adj_2191), .CO(mco_13_adj_2192), .P0(mult_10u_9u_0_pp_3_9_adj_1952), 
          .P1(mult_10u_9u_0_pp_3_10_adj_1951)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_6_2_adj_438 (.A0(VRAM_DATA_OUT[24]), .A1(VRAM_DATA_OUT[25]), 
          .A2(VRAM_DATA_OUT[25]), .A3(VRAM_DATA_OUT[26]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_13_adj_2192), .CO(mco_14_adj_2193), .P0(mult_10u_9u_0_pp_3_11_adj_1945), 
          .P1(mult_10u_9u_0_pp_3_12_adj_1944)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_6_3_adj_439 (.A0(VRAM_DATA_OUT[26]), .A1(VRAM_DATA_OUT[27]), 
          .A2(VRAM_DATA_OUT[27]), .A3(VRAM_DATA_OUT[28]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_14_adj_2193), .CO(mco_15_adj_2194), .P0(mult_10u_9u_0_pp_3_13_adj_1938), 
          .P1(mult_10u_9u_0_pp_3_14_adj_1937)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    MULT2 mult_10u_9u_0_mult_6_4_adj_440 (.A0(VRAM_DATA_OUT[28]), .A1(VRAM_DATA_OUT[29]), 
          .A2(VRAM_DATA_OUT[29]), .A3(GND_net), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_15_adj_2194), .CO(mfco_3_adj_2001), .P0(mult_10u_9u_0_pp_3_15_adj_1933), 
          .P1(mult_10u_9u_0_pp_3_16_adj_1932)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    AND2 AND2_t8_adj_441 (.A(VRAM_DATA_OUT[21]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_9_adj_2165)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(180[10:64])
    AND2 AND2_t7_adj_442 (.A(VRAM_DATA_OUT[22]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_10_adj_2166)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(182[10:65])
    AND2 AND2_t6_adj_443 (.A(VRAM_DATA_OUT[23]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_11_adj_2168)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(184[10:65])
    AND2 AND2_t5_adj_444 (.A(VRAM_DATA_OUT[24]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_12_adj_2169)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(186[10:65])
    AND2 AND2_t4_adj_445 (.A(VRAM_DATA_OUT[25]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_13_adj_2171)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(188[10:65])
    AND2 AND2_t3_adj_446 (.A(VRAM_DATA_OUT[26]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_14_adj_2172)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(190[10:65])
    AND2 AND2_t2_adj_447 (.A(VRAM_DATA_OUT[27]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_15_adj_2174)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(192[10:65])
    AND2 AND2_t1_adj_448 (.A(VRAM_DATA_OUT[28]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_16_adj_2175)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(194[10:65])
    AND2 AND2_t0_adj_449 (.A(VRAM_DATA_OUT[29]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_17_adj_2177)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(196[10:65])
    FADD2B mult_10u_9u_0_cin_lr_add_0_adj_450 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_0_adj_2178)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:100])
    AND2 AND2_t9_adj_451 (.A(BLUE_READ[0]), .B(ALPHA_READ[6]), .Z(mult_9u_9u_0_pp_3_6_adj_2195)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(165[10:63])
    AND2 AND2_t10_adj_452 (.A(BLUE_READ[0]), .B(ALPHA_READ[4]), .Z(mult_9u_9u_0_pp_2_4_adj_2196)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(163[10:64])
    AND2 AND2_t11_adj_453 (.A(BLUE_READ[0]), .B(ALPHA_READ[2]), .Z(mult_9u_9u_0_pp_1_2_adj_2197)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(161[10:64])
    AND2 AND2_t12_adj_454 (.A(BLUE_READ[0]), .B(ALPHA_READ[0]), .Z(BLUE_OUT_9__N_706[0])) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(159[10:64])
    FADD2B mult_9u_9u_0_cin_lr_add_2_adj_455 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_2_adj_2198)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_cin_lr_add_4_adj_456 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_4_adj_2199)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_cin_lr_add_6_adj_457 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_6_adj_2200)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B Cadd_mult_9u_9u_0_0_1_adj_458 (.A0(GND_net), .A1(mult_9u_9u_0_pp_0_2_adj_2202), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_1_2_adj_2197), .CI(GND_net), 
           .COUT(co_mult_9u_9u_0_0_1_adj_2201), .S1(BLUE_OUT_9__N_706[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_0_2_adj_459 (.A0(mult_9u_9u_0_pp_0_3_adj_2206), 
           .A1(mult_9u_9u_0_pp_0_4_adj_2205), .B0(mult_9u_9u_0_pp_1_3_adj_2208), 
           .B1(mult_9u_9u_0_pp_1_4_adj_2207), .CI(co_mult_9u_9u_0_0_1_adj_2201), 
           .COUT(co_mult_9u_9u_0_0_2_adj_2203), .S0(BLUE_OUT_9__N_706[3]), 
           .S1(s_mult_9u_9u_0_0_4_adj_2204)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_0_3_adj_460 (.A0(mult_9u_9u_0_pp_0_5_adj_2213), 
           .A1(mult_9u_9u_0_pp_0_6_adj_2212), .B0(mult_9u_9u_0_pp_1_5_adj_2215), 
           .B1(mult_9u_9u_0_pp_1_6_adj_2214), .CI(co_mult_9u_9u_0_0_2_adj_2203), 
           .COUT(co_mult_9u_9u_0_0_3_adj_2209), .S0(s_mult_9u_9u_0_0_5_adj_2210), 
           .S1(s_mult_9u_9u_0_0_6_adj_2211)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_0_4_adj_461 (.A0(mult_9u_9u_0_pp_0_7_adj_2220), 
           .A1(mult_9u_9u_0_pp_0_8_adj_2219), .B0(mult_9u_9u_0_pp_1_7_adj_2222), 
           .B1(mult_9u_9u_0_pp_1_8_adj_2221), .CI(co_mult_9u_9u_0_0_3_adj_2209), 
           .COUT(co_mult_9u_9u_0_0_4_adj_2216), .S0(s_mult_9u_9u_0_0_7_adj_2217), 
           .S1(s_mult_9u_9u_0_0_8_adj_2218)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_0_5_adj_462 (.A0(mult_9u_9u_0_pp_0_9_adj_2227), 
           .A1(mult_9u_9u_0_pp_0_10_adj_2226), .B0(mult_9u_9u_0_pp_1_9_adj_2229), 
           .B1(mult_9u_9u_0_pp_1_10_adj_2228), .CI(co_mult_9u_9u_0_0_4_adj_2216), 
           .COUT(co_mult_9u_9u_0_0_5_adj_2223), .S0(s_mult_9u_9u_0_0_9_adj_2224), 
           .S1(s_mult_9u_9u_0_0_10_adj_2225)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_0_6_adj_463 (.A0(GND_net), .A1(GND_net), .B0(mult_9u_9u_0_pp_1_11_adj_2234), 
           .B1(mult_9u_9u_0_pp_1_12_adj_2233), .CI(co_mult_9u_9u_0_0_5_adj_2223), 
           .COUT(co_mult_9u_9u_0_0_6_adj_2230), .S0(s_mult_9u_9u_0_0_11_adj_2231), 
           .S1(s_mult_9u_9u_0_0_12_adj_2232)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B Cadd_mult_9u_9u_0_0_7_adj_464 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_0_6_adj_2230), .S0(s_mult_9u_9u_0_0_13_adj_2235)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B Cadd_mult_9u_9u_0_1_1_adj_465 (.A0(GND_net), .A1(mult_9u_9u_0_pp_2_6_adj_2238), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_3_6_adj_2195), .CI(GND_net), 
           .COUT(co_mult_9u_9u_0_1_1_adj_2236), .S1(s_mult_9u_9u_0_1_6_adj_2237)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_1_2_adj_466 (.A0(mult_9u_9u_0_pp_2_7_adj_2243), 
           .A1(mult_9u_9u_0_pp_2_8_adj_2242), .B0(mult_9u_9u_0_pp_3_7_adj_2245), 
           .B1(mult_9u_9u_0_pp_3_8_adj_2244), .CI(co_mult_9u_9u_0_1_1_adj_2236), 
           .COUT(co_mult_9u_9u_0_1_2_adj_2239), .S0(s_mult_9u_9u_0_1_7_adj_2240), 
           .S1(s_mult_9u_9u_0_1_8_adj_2241)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_1_3_adj_467 (.A0(mult_9u_9u_0_pp_2_9_adj_2250), 
           .A1(mult_9u_9u_0_pp_2_10_adj_2249), .B0(mult_9u_9u_0_pp_3_9_adj_2252), 
           .B1(mult_9u_9u_0_pp_3_10_adj_2251), .CI(co_mult_9u_9u_0_1_2_adj_2239), 
           .COUT(co_mult_9u_9u_0_1_3_adj_2246), .S0(s_mult_9u_9u_0_1_9_adj_2247), 
           .S1(s_mult_9u_9u_0_1_10_adj_2248)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_1_4_adj_468 (.A0(mult_9u_9u_0_pp_2_11_adj_2257), 
           .A1(mult_9u_9u_0_pp_2_12_adj_2256), .B0(mult_9u_9u_0_pp_3_11_adj_2259), 
           .B1(mult_9u_9u_0_pp_3_12_adj_2258), .CI(co_mult_9u_9u_0_1_3_adj_2246), 
           .COUT(co_mult_9u_9u_0_1_4_adj_2253), .S0(s_mult_9u_9u_0_1_11_adj_2254), 
           .S1(s_mult_9u_9u_0_1_12_adj_2255)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_1_5_adj_469 (.A0(mult_9u_9u_0_pp_2_13_adj_2264), 
           .A1(mult_9u_9u_0_pp_2_14_adj_2263), .B0(mult_9u_9u_0_pp_3_13_adj_2266), 
           .B1(mult_9u_9u_0_pp_3_14_adj_2265), .CI(co_mult_9u_9u_0_1_4_adj_2253), 
           .COUT(co_mult_9u_9u_0_1_5_adj_2260), .S0(s_mult_9u_9u_0_1_13_adj_2261), 
           .S1(s_mult_9u_9u_0_1_14_adj_2262)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_1_6_adj_470 (.A0(GND_net), .A1(GND_net), .B0(mult_9u_9u_0_pp_3_15_adj_2271), 
           .B1(mult_9u_9u_0_pp_3_16_adj_2270), .CI(co_mult_9u_9u_0_1_5_adj_2260), 
           .COUT(co_mult_9u_9u_0_1_6_adj_2267), .S0(s_mult_9u_9u_0_1_15_adj_2268), 
           .S1(s_mult_9u_9u_0_1_16_adj_2269)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B Cadd_mult_9u_9u_0_1_7_adj_471 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_1_6_adj_2267), .S0(s_mult_9u_9u_0_1_17_adj_2272)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B Cadd_mult_9u_9u_0_2_1_adj_472 (.A0(GND_net), .A1(s_mult_9u_9u_0_0_4_adj_2204), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_2_4_adj_2196), .CI(GND_net), 
           .COUT(co_mult_9u_9u_0_2_1_adj_2273), .S1(BLUE_OUT_9__N_706[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_2_adj_473 (.A0(s_mult_9u_9u_0_0_5_adj_2210), 
           .A1(s_mult_9u_9u_0_0_6_adj_2211), .B0(mult_9u_9u_0_pp_2_5_adj_2275), 
           .B1(s_mult_9u_9u_0_1_6_adj_2237), .CI(co_mult_9u_9u_0_2_1_adj_2273), 
           .COUT(co_mult_9u_9u_0_2_2_adj_2274), .S0(BLUE_OUT_9__N_706[5]), 
           .S1(BLUE_OUT_9__N_706[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_3_adj_474 (.A0(s_mult_9u_9u_0_0_7_adj_2217), 
           .A1(s_mult_9u_9u_0_0_8_adj_2218), .B0(s_mult_9u_9u_0_1_7_adj_2240), 
           .B1(s_mult_9u_9u_0_1_8_adj_2241), .CI(co_mult_9u_9u_0_2_2_adj_2274), 
           .COUT(co_mult_9u_9u_0_2_3_adj_2276), .S0(BLUE_OUT_9__N_706[7]), 
           .S1(s_mult_9u_9u_0_2_8_adj_2277)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_4_adj_475 (.A0(s_mult_9u_9u_0_0_9_adj_2224), 
           .A1(s_mult_9u_9u_0_0_10_adj_2225), .B0(s_mult_9u_9u_0_1_9_adj_2247), 
           .B1(s_mult_9u_9u_0_1_10_adj_2248), .CI(co_mult_9u_9u_0_2_3_adj_2276), 
           .COUT(co_mult_9u_9u_0_2_4_adj_2278), .S0(s_mult_9u_9u_0_2_9_adj_2279), 
           .S1(s_mult_9u_9u_0_2_10_adj_2280)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_5_adj_476 (.A0(s_mult_9u_9u_0_0_11_adj_2231), 
           .A1(s_mult_9u_9u_0_0_12_adj_2232), .B0(s_mult_9u_9u_0_1_11_adj_2254), 
           .B1(s_mult_9u_9u_0_1_12_adj_2255), .CI(co_mult_9u_9u_0_2_4_adj_2278), 
           .COUT(co_mult_9u_9u_0_2_5_adj_2281), .S0(s_mult_9u_9u_0_2_11_adj_2282), 
           .S1(s_mult_9u_9u_0_2_12_adj_2283)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_6_adj_477 (.A0(s_mult_9u_9u_0_0_13_adj_2235), 
           .A1(GND_net), .B0(s_mult_9u_9u_0_1_13_adj_2261), .B1(s_mult_9u_9u_0_1_14_adj_2262), 
           .CI(co_mult_9u_9u_0_2_5_adj_2281), .COUT(co_mult_9u_9u_0_2_6_adj_2284), 
           .S0(s_mult_9u_9u_0_2_13_adj_2285), .S1(s_mult_9u_9u_0_2_14_adj_2286)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_7_adj_478 (.A0(GND_net), .A1(GND_net), .B0(s_mult_9u_9u_0_1_15_adj_2268), 
           .B1(s_mult_9u_9u_0_1_16_adj_2269), .CI(co_mult_9u_9u_0_2_6_adj_2284), 
           .COUT(co_mult_9u_9u_0_2_7_adj_2287), .S0(s_mult_9u_9u_0_2_15_adj_2288), 
           .S1(s_mult_9u_9u_0_2_16_adj_2289)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B mult_9u_9u_0_add_2_8_adj_479 (.A0(GND_net), .A1(GND_net), .B0(s_mult_9u_9u_0_1_17_adj_2272), 
           .B1(GND_net), .CI(co_mult_9u_9u_0_2_7_adj_2287), .S0(s_mult_9u_9u_0_2_17_adj_2290)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B Cadd_t_mult_9u_9u_0_3_1_adj_480 (.A0(GND_net), .A1(s_mult_9u_9u_0_2_8_adj_2277), 
           .B0(GND_net), .B1(mult_9u_9u_0_pp_4_8_adj_1882), .CI(GND_net), 
           .COUT(co_t_mult_9u_9u_0_3_1_adj_2291), .S1(BLUE_OUT_9__N_706[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B t_mult_9u_9u_0_add_3_2_adj_481 (.A0(s_mult_9u_9u_0_2_9_adj_2279), 
           .A1(s_mult_9u_9u_0_2_10_adj_2280), .B0(mult_9u_9u_0_pp_4_9_adj_2292), 
           .B1(mult_9u_9u_0_pp_4_10_adj_2293), .CI(co_t_mult_9u_9u_0_3_1_adj_2291), 
           .COUT(co_t_mult_9u_9u_0_3_2_adj_2294), .S0(BLUE_OUT_9__N_706[9]), 
           .S1(BLUE_OUT_9__N_706[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B t_mult_9u_9u_0_add_3_3_adj_482 (.A0(s_mult_9u_9u_0_2_11_adj_2282), 
           .A1(s_mult_9u_9u_0_2_12_adj_2283), .B0(mult_9u_9u_0_pp_4_11_adj_2295), 
           .B1(mult_9u_9u_0_pp_4_12_adj_2296), .CI(co_t_mult_9u_9u_0_3_2_adj_2294), 
           .COUT(co_t_mult_9u_9u_0_3_3_adj_2297), .S0(BLUE_OUT_9__N_706[11]), 
           .S1(BLUE_OUT_9__N_706[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B t_mult_9u_9u_0_add_3_4_adj_483 (.A0(s_mult_9u_9u_0_2_13_adj_2285), 
           .A1(s_mult_9u_9u_0_2_14_adj_2286), .B0(mult_9u_9u_0_pp_4_13_adj_2298), 
           .B1(mult_9u_9u_0_pp_4_14_adj_2299), .CI(co_t_mult_9u_9u_0_3_3_adj_2297), 
           .COUT(co_t_mult_9u_9u_0_3_4_adj_2300), .S0(BLUE_OUT_9__N_706[13]), 
           .S1(BLUE_OUT_9__N_706[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B t_mult_9u_9u_0_add_3_5_adj_484 (.A0(s_mult_9u_9u_0_2_15_adj_2288), 
           .A1(s_mult_9u_9u_0_2_16_adj_2289), .B0(mult_9u_9u_0_pp_4_15_adj_2301), 
           .B1(mult_9u_9u_0_pp_4_16_adj_2302), .CI(co_t_mult_9u_9u_0_3_4_adj_2300), 
           .COUT(co_t_mult_9u_9u_0_3_5_adj_2303), .S0(BLUE_OUT_9__N_706[15]), 
           .S1(BLUE_OUT_9__N_706[16])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    FADD2B t_mult_9u_9u_0_add_3_6_adj_485 (.A0(s_mult_9u_9u_0_2_17_adj_2290), 
           .A1(GND_net), .B0(GND_net), .B1(GND_net), .CI(co_t_mult_9u_9u_0_3_5_adj_2303), 
           .S0(BLUE_OUT_9__N_706[17])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_0_0_adj_486 (.A0(BLUE_READ[0]), .A1(BLUE_READ[1]), 
          .A2(BLUE_READ[1]), .A3(BLUE_READ[2]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), 
          .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), .CI(mult_9u_9u_0_cin_lr_0_adj_2304), 
          .CO(mco_adj_2305), .P0(BLUE_OUT_9__N_706[1]), .P1(mult_9u_9u_0_pp_0_2_adj_2202)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_0_1_adj_487 (.A0(BLUE_READ[2]), .A1(BLUE_READ[3]), 
          .A2(BLUE_READ[3]), .A3(BLUE_READ[4]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), 
          .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), .CI(mco_adj_2305), .CO(mco_1_adj_2306), 
          .P0(mult_9u_9u_0_pp_0_3_adj_2206), .P1(mult_9u_9u_0_pp_0_4_adj_2205)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_0_2_adj_488 (.A0(BLUE_READ[4]), .A1(BLUE_READ[5]), 
          .A2(BLUE_READ[5]), .A3(BLUE_READ[6]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), 
          .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), .CI(mco_1_adj_2306), 
          .CO(mco_2_adj_2307), .P0(mult_9u_9u_0_pp_0_5_adj_2213), .P1(mult_9u_9u_0_pp_0_6_adj_2212)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_0_3_adj_489 (.A0(BLUE_READ[6]), .A1(BLUE_READ[7]), 
          .A2(BLUE_READ[7]), .A3(BLUE_READ[8]), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), 
          .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), .CI(mco_2_adj_2307), 
          .CO(mco_3_adj_2308), .P0(mult_9u_9u_0_pp_0_7_adj_2220), .P1(mult_9u_9u_0_pp_0_8_adj_2219)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_0_4_adj_490 (.A0(BLUE_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[1]), .B1(ALPHA_READ[0]), 
          .B2(ALPHA_READ[1]), .B3(ALPHA_READ[0]), .CI(mco_3_adj_2308), 
          .P0(mult_9u_9u_0_pp_0_9_adj_2227), .P1(mult_9u_9u_0_pp_0_10_adj_2226)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_2_0_adj_491 (.A0(BLUE_READ[0]), .A1(BLUE_READ[1]), 
          .A2(BLUE_READ[1]), .A3(BLUE_READ[2]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), 
          .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), .CI(mult_9u_9u_0_cin_lr_2_adj_2198), 
          .CO(mco_4_adj_2309), .P0(mult_9u_9u_0_pp_1_3_adj_2208), .P1(mult_9u_9u_0_pp_1_4_adj_2207)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_2_1_adj_492 (.A0(BLUE_READ[2]), .A1(BLUE_READ[3]), 
          .A2(BLUE_READ[3]), .A3(BLUE_READ[4]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), 
          .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), .CI(mco_4_adj_2309), 
          .CO(mco_5_adj_2310), .P0(mult_9u_9u_0_pp_1_5_adj_2215), .P1(mult_9u_9u_0_pp_1_6_adj_2214)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_2_2_adj_493 (.A0(BLUE_READ[4]), .A1(BLUE_READ[5]), 
          .A2(BLUE_READ[5]), .A3(BLUE_READ[6]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), 
          .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), .CI(mco_5_adj_2310), 
          .CO(mco_6_adj_2311), .P0(mult_9u_9u_0_pp_1_7_adj_2222), .P1(mult_9u_9u_0_pp_1_8_adj_2221)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_2_3_adj_494 (.A0(BLUE_READ[6]), .A1(BLUE_READ[7]), 
          .A2(BLUE_READ[7]), .A3(BLUE_READ[8]), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), 
          .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), .CI(mco_6_adj_2311), 
          .CO(mco_7_adj_2312), .P0(mult_9u_9u_0_pp_1_9_adj_2229), .P1(mult_9u_9u_0_pp_1_10_adj_2228)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_2_4_adj_495 (.A0(BLUE_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[3]), .B1(ALPHA_READ[2]), 
          .B2(ALPHA_READ[3]), .B3(ALPHA_READ[2]), .CI(mco_7_adj_2312), 
          .P0(mult_9u_9u_0_pp_1_11_adj_2234), .P1(mult_9u_9u_0_pp_1_12_adj_2233)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_4_0_adj_496 (.A0(BLUE_READ[0]), .A1(BLUE_READ[1]), 
          .A2(BLUE_READ[1]), .A3(BLUE_READ[2]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), 
          .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), .CI(mult_9u_9u_0_cin_lr_4_adj_2199), 
          .CO(mco_8_adj_2313), .P0(mult_9u_9u_0_pp_2_5_adj_2275), .P1(mult_9u_9u_0_pp_2_6_adj_2238)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_4_1_adj_497 (.A0(BLUE_READ[2]), .A1(BLUE_READ[3]), 
          .A2(BLUE_READ[3]), .A3(BLUE_READ[4]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), 
          .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), .CI(mco_8_adj_2313), 
          .CO(mco_9_adj_2314), .P0(mult_9u_9u_0_pp_2_7_adj_2243), .P1(mult_9u_9u_0_pp_2_8_adj_2242)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_4_2_adj_498 (.A0(BLUE_READ[4]), .A1(BLUE_READ[5]), 
          .A2(BLUE_READ[5]), .A3(BLUE_READ[6]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), 
          .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), .CI(mco_9_adj_2314), 
          .CO(mco_10_adj_2315), .P0(mult_9u_9u_0_pp_2_9_adj_2250), .P1(mult_9u_9u_0_pp_2_10_adj_2249)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_4_3_adj_499 (.A0(BLUE_READ[6]), .A1(BLUE_READ[7]), 
          .A2(BLUE_READ[7]), .A3(BLUE_READ[8]), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), 
          .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), .CI(mco_10_adj_2315), 
          .CO(mco_11_adj_2316), .P0(mult_9u_9u_0_pp_2_11_adj_2257), .P1(mult_9u_9u_0_pp_2_12_adj_2256)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_4_4_adj_500 (.A0(BLUE_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[5]), .B1(ALPHA_READ[4]), 
          .B2(ALPHA_READ[5]), .B3(ALPHA_READ[4]), .CI(mco_11_adj_2316), 
          .P0(mult_9u_9u_0_pp_2_13_adj_2264), .P1(mult_9u_9u_0_pp_2_14_adj_2263)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_6_0_adj_501 (.A0(BLUE_READ[0]), .A1(BLUE_READ[1]), 
          .A2(BLUE_READ[1]), .A3(BLUE_READ[2]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), 
          .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), .CI(mult_9u_9u_0_cin_lr_6_adj_2200), 
          .CO(mco_12_adj_2317), .P0(mult_9u_9u_0_pp_3_7_adj_2245), .P1(mult_9u_9u_0_pp_3_8_adj_2244)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_6_1_adj_502 (.A0(BLUE_READ[2]), .A1(BLUE_READ[3]), 
          .A2(BLUE_READ[3]), .A3(BLUE_READ[4]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), 
          .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), .CI(mco_12_adj_2317), 
          .CO(mco_13_adj_2318), .P0(mult_9u_9u_0_pp_3_9_adj_2252), .P1(mult_9u_9u_0_pp_3_10_adj_2251)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_6_2_adj_503 (.A0(BLUE_READ[4]), .A1(BLUE_READ[5]), 
          .A2(BLUE_READ[5]), .A3(BLUE_READ[6]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), 
          .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), .CI(mco_13_adj_2318), 
          .CO(mco_14_adj_2319), .P0(mult_9u_9u_0_pp_3_11_adj_2259), .P1(mult_9u_9u_0_pp_3_12_adj_2258)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_6_3_adj_504 (.A0(BLUE_READ[6]), .A1(BLUE_READ[7]), 
          .A2(BLUE_READ[7]), .A3(BLUE_READ[8]), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), 
          .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), .CI(mco_14_adj_2319), 
          .CO(mco_15_adj_2320), .P0(mult_9u_9u_0_pp_3_13_adj_2266), .P1(mult_9u_9u_0_pp_3_14_adj_2265)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    MULT2 mult_9u_9u_0_mult_6_4_adj_505 (.A0(BLUE_READ[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(ALPHA_READ[7]), .B1(ALPHA_READ[6]), 
          .B2(ALPHA_READ[7]), .B3(ALPHA_READ[6]), .CI(mco_15_adj_2320), 
          .P0(mult_9u_9u_0_pp_3_15_adj_2271), .P1(mult_9u_9u_0_pp_3_16_adj_2270)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    AND2 AND2_t7_adj_506 (.A(BLUE_READ[1]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_9_adj_2292)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(169[10:63])
    AND2 AND2_t6_adj_507 (.A(BLUE_READ[2]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_10_adj_2293)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(171[10:64])
    AND2 AND2_t5_adj_508 (.A(BLUE_READ[3]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_11_adj_2295)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(173[10:64])
    AND2 AND2_t4_adj_509 (.A(BLUE_READ[4]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_12_adj_2296)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(175[10:64])
    AND2 AND2_t3_adj_510 (.A(BLUE_READ[5]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_13_adj_2298)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(177[10:64])
    AND2 AND2_t2_adj_511 (.A(BLUE_READ[6]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_14_adj_2299)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(179[10:64])
    AND2 AND2_t1_adj_512 (.A(BLUE_READ[7]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_15_adj_2301)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(181[10:64])
    AND2 AND2_t0_adj_513 (.A(BLUE_READ[8]), .B(ALPHA_READ[8]), .Z(mult_9u_9u_0_pp_4_16_adj_2302)) /* synthesis syn_instantiated=1 */ ;   // mult_9u_9u.v(183[10:64])
    FADD2B mult_9u_9u_0_cin_lr_add_0_adj_514 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_9u_9u_0_cin_lr_0_adj_2304)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[128:148])
    LUT4 i31_2_lut (.A(BUS_transferState[1]), .B(BUS_transferState[0]), 
         .Z(n17)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i31_2_lut.init = 16'h6666;
    LUT4 i12367_3_lut (.A(n3974), .B(n3990), .C(currSprite[4]), .Z(n16029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12367_3_lut.init = 16'hcaca;
    LUT4 state_7__I_0_i13_2_lut_rep_439 (.A(state[6]), .B(state[7]), .Z(n17447)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam state_7__I_0_i13_2_lut_rep_439.init = 16'heeee;
    PFUMX i12571 (.BLUT(n16231), .ALUT(n16232), .C0(n17334), .Z(Sprite_readData2_15__N_476[0]));
    LUT4 i12366_3_lut (.A(n3939), .B(n3955), .C(currSprite[4]), .Z(n16028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12366_3_lut.init = 16'hcaca;
    LUT4 i12364_3_lut (.A(n4078), .B(n4094), .C(currSprite[4]), .Z(n16026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12364_3_lut.init = 16'hcaca;
    PFUMX i12574 (.BLUT(n16234), .ALUT(n16235), .C0(n17334), .Z(Sprite_readData2_15__N_476[1]));
    LUT4 i1_3_lut_3_lut_4_lut (.A(state[6]), .B(state[7]), .C(\state[1] ), 
         .D(\state[0] ), .Z(n5_adj_2321)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i1_3_lut_3_lut_4_lut.init = 16'heefe;
    LUT4 state_7__I_0_772_i12_2_lut_rep_440 (.A(state[4]), .B(state[5]), 
         .Z(n17448)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(365[10:23])
    defparam state_7__I_0_772_i12_2_lut_rep_440.init = 16'heeee;
    CCU2D add_10518_9 (.A0(n16[7]), .B0(\Sprite_readAddr_13__N_752[7] ), 
          .C0(GND_net), .D0(GND_net), .A1(n16[8]), .B1(\Sprite_readAddr_13__N_752[8] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14122), .COUT(n14123), .S0(Sprite_readAddr[7]), 
          .S1(Sprite_readAddr[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_9.INIT0 = 16'h5666;
    defparam add_10518_9.INIT1 = 16'h5666;
    defparam add_10518_9.INJECT1_0 = "NO";
    defparam add_10518_9.INJECT1_1 = "NO";
    CCU2D add_10518_7 (.A0(n16[5]), .B0(\Sprite_readAddr_13__N_752[5] ), 
          .C0(GND_net), .D0(GND_net), .A1(n16[6]), .B1(\Sprite_readAddr_13__N_752[6] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14121), .COUT(n14122), .S0(Sprite_readAddr[5]), 
          .S1(Sprite_readAddr[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_7.INIT0 = 16'h5666;
    defparam add_10518_7.INIT1 = 16'h5666;
    defparam add_10518_7.INJECT1_0 = "NO";
    defparam add_10518_7.INJECT1_1 = "NO";
    LUT4 i12363_3_lut (.A(n4043), .B(n4059), .C(currSprite[4]), .Z(n16025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12363_3_lut.init = 16'hcaca;
    CCU2D add_10518_5 (.A0(n16[3]), .B0(\Sprite_readAddr_13__N_752[3] ), 
          .C0(GND_net), .D0(GND_net), .A1(n16[4]), .B1(\Sprite_readAddr_13__N_752[4] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14120), .COUT(n14121), .S0(Sprite_readAddr[3]), 
          .S1(Sprite_readAddr[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_5.INIT0 = 16'h5666;
    defparam add_10518_5.INIT1 = 16'h5666;
    defparam add_10518_5.INJECT1_0 = "NO";
    defparam add_10518_5.INJECT1_1 = "NO";
    CCU2D add_10518_3 (.A0(n16[1]), .B0(\Sprite_readAddr_13__N_752[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(n16[2]), .B1(\Sprite_readAddr_13__N_752[2] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14119), .COUT(n14120), .S0(Sprite_readAddr[1]), 
          .S1(Sprite_readAddr[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_3.INIT0 = 16'h5666;
    defparam add_10518_3.INIT1 = 16'h5666;
    defparam add_10518_3.INJECT1_0 = "NO";
    defparam add_10518_3.INJECT1_1 = "NO";
    LUT4 state_7__I_0_764_i14_2_lut_rep_397_3_lut_4_lut (.A(state[4]), .B(state[5]), 
         .C(state[7]), .D(state[6]), .Z(n17405)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(365[10:23])
    defparam state_7__I_0_764_i14_2_lut_rep_397_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_515 (.A(state[4]), .B(state[5]), .C(n17275), 
         .D(\state[0] ), .Z(n15420)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(365[10:23])
    defparam i1_3_lut_4_lut_adj_515.init = 16'h0100;
    LUT4 i1_4_lut_adj_516 (.A(BUS_transferState[1]), .B(GR_WR_CLK), .C(BUS_transferState[0]), 
         .D(BUS_transferState[2]), .Z(GR_WR_CLK_N_1081)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A !(B+!((D)+!C)))) */ ;
    defparam i1_4_lut_adj_516.init = 16'h4cd4;
    LUT4 state_7__I_0_772_i9_2_lut_rep_441 (.A(\state[0] ), .B(\state[1] ), 
         .Z(n17449)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(365[10:23])
    defparam state_7__I_0_772_i9_2_lut_rep_441.init = 16'heeee;
    PFUMX i12577 (.BLUT(n16237), .ALUT(n16238), .C0(n17334), .Z(Sprite_readData2_15__N_476[2]));
    LUT4 i2_3_lut_4_lut_adj_517 (.A(\state[0] ), .B(\state[1] ), .C(state[2]), 
         .D(\state[3] ), .Z(n15508)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(365[10:23])
    defparam i2_3_lut_4_lut_adj_517.init = 16'hffef;
    LUT4 state_7__I_0_i10_2_lut_rep_442 (.A(state[2]), .B(\state[3] ), .Z(n17450)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam state_7__I_0_i10_2_lut_rep_442.init = 16'heeee;
    LUT4 i1_2_lut_rep_395_3_lut_4_lut (.A(state[2]), .B(\state[3] ), .C(\state[1] ), 
         .D(\state[0] ), .Z(n17403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i1_2_lut_rep_395_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12361_3_lut (.A(n4081), .B(n4097), .C(currSprite[4]), .Z(n16023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12361_3_lut.init = 16'hcaca;
    LUT4 i12360_3_lut (.A(n4046), .B(n4062), .C(currSprite[4]), .Z(n16022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12360_3_lut.init = 16'hcaca;
    CCU2D add_10518_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(SpriteRead_xInSprite[0]), .B1(n3855[0]), .C1(\Sprite_readAddr_13__N_752[0] ), 
          .D1(GND_net), .COUT(n14119), .S1(Sprite_readAddr[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_10518_1.INIT0 = 16'hF000;
    defparam add_10518_1.INIT1 = 16'h9696;
    defparam add_10518_1.INJECT1_0 = "NO";
    defparam add_10518_1.INJECT1_1 = "NO";
    CCU2D BLUE_OUT_9__I_0_10 (.A0(BLUE_OUT_9__N_687[8]), .B0(BLUE_OUT_9__N_706[8]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[9]), .B1(BLUE_OUT_9__N_706[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14051), .COUT(n14052), .S1(BLUE_OUT[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_10.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_10.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_10.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_10.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_396_3_lut (.A(state[2]), .B(\state[3] ), .C(\state[1] ), 
         .Z(n17404)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i1_2_lut_rep_396_3_lut.init = 16'hfefe;
    LUT4 i12358_3_lut (.A(n3969), .B(n3985), .C(currSprite[4]), .Z(n16020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12358_3_lut.init = 16'hcaca;
    PFUMX i13398 (.BLUT(n17256), .ALUT(n17255), .C0(\state[0] ), .Z(n17257));
    LUT4 i2_2_lut_rep_359_3_lut_4_lut (.A(state[2]), .B(\state[3] ), .C(\state[0] ), 
         .D(\state[1] ), .Z(n17367)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i2_2_lut_rep_359_3_lut_4_lut.init = 16'hffef;
    PFUMX i12580 (.BLUT(n16240), .ALUT(n16241), .C0(n17334), .Z(Sprite_readData2_15__N_476[3]));
    LUT4 i12357_3_lut (.A(n3934), .B(n3950), .C(currSprite[4]), .Z(n16019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12357_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_443 (.A(state[5]), .B(\state[1] ), .C(state[6]), 
         .Z(n17451)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam i2_3_lut_rep_443.init = 16'h8080;
    CCU2D BLUE_OUT_9__I_0_8 (.A0(BLUE_OUT_9__N_687[6]), .B0(BLUE_OUT_9__N_706[6]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[7]), .B1(BLUE_OUT_9__N_706[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14050), .COUT(n14051));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_8.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_8.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_8.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_8.INJECT1_1 = "NO";
    PFUMX i12583 (.BLUT(n16243), .ALUT(n16244), .C0(n17334), .Z(Sprite_readData2_15__N_476[4]));
    PFUMX i12586 (.BLUT(n16246), .ALUT(n16247), .C0(n17334), .Z(Sprite_readData2_15__N_476[5]));
    CCU2D BLUE_OUT_9__I_0_6 (.A0(BLUE_OUT_9__N_687[4]), .B0(BLUE_OUT_9__N_706[4]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[5]), .B1(BLUE_OUT_9__N_706[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14049), .COUT(n14050));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_6.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_6.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_6.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_6.INJECT1_1 = "NO";
    CCU2D BLUE_OUT_9__I_0_4 (.A0(BLUE_OUT_9__N_687[2]), .B0(BLUE_OUT_9__N_706[2]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[3]), .B1(BLUE_OUT_9__N_706[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14048), .COUT(n14049));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_4.INIT0 = 16'h5666;
    defparam BLUE_OUT_9__I_0_4.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_4.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_4.INJECT1_1 = "NO";
    PFUMX i12592 (.BLUT(n16251), .ALUT(n16252), .C0(n17342), .Z(n16254));
    LUT4 i12355_3_lut (.A(n3971), .B(n3987), .C(currSprite[4]), .Z(n16017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12355_3_lut.init = 16'hcaca;
    PFUMX i12596 (.BLUT(n16256), .ALUT(n16257), .C0(n17334), .Z(Sprite_readData2_15__N_476[6]));
    LUT4 i12354_3_lut (.A(n3936), .B(n3952), .C(currSprite[4]), .Z(n16016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12354_3_lut.init = 16'hcaca;
    LUT4 LED_c_bdd_2_lut_13367_3_lut (.A(n17175), .B(n2539), .C(n15352), 
         .Z(LOGIC_CLOCK_enable_51)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam LED_c_bdd_2_lut_13367_3_lut.init = 16'h2020;
    LUT4 i12352_3_lut (.A(n3963), .B(n3979), .C(currSprite[4]), .Z(n16014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12352_3_lut.init = 16'hcaca;
    PFUMX i12599 (.BLUT(n16259), .ALUT(n16260), .C0(n17334), .Z(Sprite_readData2_15__N_476[7]));
    LUT4 i12351_3_lut (.A(n3928), .B(n3944), .C(currSprite[4]), .Z(n16013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12351_3_lut.init = 16'hcaca;
    PFUMX i12602 (.BLUT(n16262), .ALUT(n16263), .C0(n17334), .Z(Sprite_readData2_15__N_476[8]));
    LUT4 i12349_3_lut (.A(n3976), .B(n3992), .C(currSprite[4]), .Z(n16011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12349_3_lut.init = 16'hcaca;
    LUT4 i12348_3_lut (.A(n3941), .B(n3957), .C(currSprite[4]), .Z(n16010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12348_3_lut.init = 16'hcaca;
    PFUMX i12107 (.BLUT(n15767), .ALUT(n15768), .C0(n17334), .Z(Sprite_readData2_15__N_524[7]));
    LUT4 i12346_3_lut (.A(n3964), .B(n3980), .C(currSprite[4]), .Z(n16008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12346_3_lut.init = 16'hcaca;
    LUT4 i12345_3_lut (.A(n3929), .B(n3945), .C(currSprite[4]), .Z(n16007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12345_3_lut.init = 16'hcaca;
    LUT4 i6680_2_lut_rep_446 (.A(BUS_transferState[0]), .B(BUS_transferState[1]), 
         .Z(n17454)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6680_2_lut_rep_446.init = 16'h8888;
    PFUMX i12605 (.BLUT(n16265), .ALUT(n16266), .C0(n17334), .Z(Sprite_readData2_15__N_492[0]));
    LUT4 i1_2_lut_4_lut_adj_518 (.A(n17287), .B(n17428), .C(n17286), .D(n17306), 
         .Z(n15448)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[4] 608[11])
    defparam i1_2_lut_4_lut_adj_518.init = 16'h003a;
    LUT4 i12343_3_lut (.A(n4080), .B(n4096), .C(currSprite[4]), .Z(n16005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12343_3_lut.init = 16'hcaca;
    CCU2D BLUE_OUT_9__I_0_2 (.A0(BLUE_OUT_9__N_687[0]), .B0(BLUE_OUT_9__N_706[0]), 
          .C0(GND_net), .D0(GND_net), .A1(BLUE_OUT_9__N_687[1]), .B1(BLUE_OUT_9__N_706[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n14048));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[36:101])
    defparam BLUE_OUT_9__I_0_2.INIT0 = 16'h7000;
    defparam BLUE_OUT_9__I_0_2.INIT1 = 16'h5666;
    defparam BLUE_OUT_9__I_0_2.INJECT1_0 = "NO";
    defparam BLUE_OUT_9__I_0_2.INJECT1_1 = "NO";
    PFUMX i12110 (.BLUT(n15770), .ALUT(n15771), .C0(n17334), .Z(Sprite_readData2_15__N_524[8]));
    LUT4 i12342_3_lut (.A(n4045), .B(n4061), .C(currSprite[4]), .Z(n16004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12342_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut (.A(BUS_transferState[0]), .B(BUS_transferState[1]), 
         .C(BUS_transferState[2]), .Z(n5113)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i12340_3_lut (.A(n3965), .B(n3981), .C(currSprite[4]), .Z(n16002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12340_3_lut.init = 16'hcaca;
    CCU2D sub_47_add_2_9 (.A0(xPre[7]), .B0(currSprite_pos[7]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14113), .S0(SpriteRead_xInSprite[7]), .S1(SpriteRead_xValid_N_1166));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(273[43:57])
    defparam sub_47_add_2_9.INIT0 = 16'h5999;
    defparam sub_47_add_2_9.INIT1 = 16'h0000;
    defparam sub_47_add_2_9.INJECT1_0 = "NO";
    defparam sub_47_add_2_9.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_20 (.A0(GREEN_OUT_9__N_650[18]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14047), .S0(GREEN_OUT[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_20.INIT0 = 16'h5aaa;
    defparam GREEN_OUT_9__I_0_20.INIT1 = 16'h0000;
    defparam GREEN_OUT_9__I_0_20.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_20.INJECT1_1 = "NO";
    LUT4 i2451_2_lut (.A(BUS_transferState[2]), .B(BUS_transferState[1]), 
         .Z(BUS_transferState_3__N_930[2])) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(583[5] 607[12])
    defparam i2451_2_lut.init = 16'heeee;
    CCU2D add_10513_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13]_adj_7 ), .D0(n18266), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14]_adj_3 ), 
          .D1(n18262), .CIN(n13998), .COUT(n13999));
    defparam add_10513_7.INIT0 = 16'h00ce;
    defparam add_10513_7.INIT1 = 16'h00ce;
    defparam add_10513_7.INJECT1_0 = "NO";
    defparam add_10513_7.INJECT1_1 = "NO";
    PFUMX i12611 (.BLUT(n16270), .ALUT(n16271), .C0(n17342), .Z(n16273));
    CCU2D sub_47_add_2_7 (.A0(xPre[5]), .B0(currSprite_pos[5]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[6]), .B1(currSprite_pos[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14112), .COUT(n14113), .S0(SpriteRead_xInSprite[5]), 
          .S1(SpriteRead_xInSprite[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(273[43:57])
    defparam sub_47_add_2_7.INIT0 = 16'h5999;
    defparam sub_47_add_2_7.INIT1 = 16'h5999;
    defparam sub_47_add_2_7.INJECT1_0 = "NO";
    defparam sub_47_add_2_7.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_18 (.A0(GREEN_OUT_9__N_650[16]), .B0(GREEN_OUT_9__N_669[16]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[17]), .B1(GREEN_OUT_9__N_669[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14046), .COUT(n14047), .S0(GREEN_OUT[7]), 
          .S1(GREEN_OUT[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_18.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_18.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_18.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_18.INJECT1_1 = "NO";
    LUT4 i12339_3_lut (.A(n3930), .B(n3946), .C(currSprite[4]), .Z(n16001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12339_3_lut.init = 16'hcaca;
    LUT4 i12337_3_lut (.A(n3966), .B(n3982), .C(currSprite[4]), .Z(n15999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12337_3_lut.init = 16'hcaca;
    LUT4 i12336_3_lut (.A(n3931), .B(n3947), .C(currSprite[4]), .Z(n15998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12336_3_lut.init = 16'hcaca;
    PFUMX i12615 (.BLUT(n16275), .ALUT(n16276), .C0(n17334), .Z(Sprite_readData2_15__N_492[1]));
    LUT4 i12334_3_lut (.A(n3967), .B(n3983), .C(currSprite[4]), .Z(n15996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12334_3_lut.init = 16'hcaca;
    LUT4 i12038_3_lut (.A(\state[1] ), .B(\state[3] ), .C(\state[0] ), 
         .Z(n15699)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i12038_3_lut.init = 16'hfefe;
    CCU2D sub_47_add_2_5 (.A0(xPre[3]), .B0(currSprite_pos[3]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[4]), .B1(currSprite_pos[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14111), .COUT(n14112), .S0(SpriteRead_xInSprite[3]), 
          .S1(SpriteRead_xInSprite[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(273[43:57])
    defparam sub_47_add_2_5.INIT0 = 16'h5999;
    defparam sub_47_add_2_5.INIT1 = 16'h5999;
    defparam sub_47_add_2_5.INJECT1_0 = "NO";
    defparam sub_47_add_2_5.INJECT1_1 = "NO";
    LUT4 i12333_3_lut (.A(n3932), .B(n3948), .C(currSprite[4]), .Z(n15995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12333_3_lut.init = 16'hcaca;
    PFUMX i12618 (.BLUT(n16278), .ALUT(n16279), .C0(n17334), .Z(Sprite_readData2_15__N_492[2]));
    AND2 AND2_t10_adj_519 (.A(VRAM_DATA_OUT[0]), .B(RED_OUT_9__N_768[6]), 
         .Z(mult_10u_9u_0_pp_3_6_adj_2322)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(176[10:65])
    AND2 AND2_t11_adj_520 (.A(VRAM_DATA_OUT[0]), .B(RED_OUT_9__N_768[4]), 
         .Z(mult_10u_9u_0_pp_2_4_adj_2323)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(174[10:65])
    AND2 AND2_t12_adj_521 (.A(VRAM_DATA_OUT[0]), .B(RED_OUT_9__N_768[2]), 
         .Z(mult_10u_9u_0_pp_1_2_adj_2324)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(172[10:65])
    AND2 AND2_t13_adj_522 (.A(VRAM_DATA_OUT[0]), .B(RED_OUT_9__N_768[0]), 
         .Z(RED_OUT_9__N_613[0])) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(170[10:65])
    FADD2B mult_10u_9u_0_Cadd_0_5_adj_523 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_adj_2326), .S0(mult_10u_9u_0_pp_0_11_adj_2325)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_cin_lr_add_2_adj_524 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_2_adj_2327)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_Cadd_2_5_adj_525 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1_adj_2329), .S0(mult_10u_9u_0_pp_1_13_adj_2328)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_cin_lr_add_4_adj_526 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_4_adj_2330)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_Cadd_4_5_adj_527 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2_adj_2332), .S0(mult_10u_9u_0_pp_2_15_adj_2331)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_cin_lr_add_6_adj_528 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_6_adj_2333)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_Cadd_6_5_adj_529 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3_adj_2335), .S0(mult_10u_9u_0_pp_3_17_adj_2334)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B Cadd_mult_10u_9u_0_0_1_adj_530 (.A0(GND_net), .A1(mult_10u_9u_0_pp_0_2_adj_2337), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_1_2_adj_2324), .CI(GND_net), 
           .COUT(co_mult_10u_9u_0_0_1_adj_2336), .S1(RED_OUT_9__N_613[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_0_2_adj_531 (.A0(mult_10u_9u_0_pp_0_3_adj_2341), 
           .A1(mult_10u_9u_0_pp_0_4_adj_2340), .B0(mult_10u_9u_0_pp_1_3_adj_2343), 
           .B1(mult_10u_9u_0_pp_1_4_adj_2342), .CI(co_mult_10u_9u_0_0_1_adj_2336), 
           .COUT(co_mult_10u_9u_0_0_2_adj_2338), .S0(RED_OUT_9__N_613[3]), 
           .S1(s_mult_10u_9u_0_0_4_adj_2339)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_0_3_adj_532 (.A0(mult_10u_9u_0_pp_0_5_adj_2348), 
           .A1(mult_10u_9u_0_pp_0_6_adj_2347), .B0(mult_10u_9u_0_pp_1_5_adj_2350), 
           .B1(mult_10u_9u_0_pp_1_6_adj_2349), .CI(co_mult_10u_9u_0_0_2_adj_2338), 
           .COUT(co_mult_10u_9u_0_0_3_adj_2344), .S0(s_mult_10u_9u_0_0_5_adj_2345), 
           .S1(s_mult_10u_9u_0_0_6_adj_2346)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_0_4_adj_533 (.A0(mult_10u_9u_0_pp_0_7_adj_2355), 
           .A1(mult_10u_9u_0_pp_0_8_adj_2354), .B0(mult_10u_9u_0_pp_1_7_adj_2357), 
           .B1(mult_10u_9u_0_pp_1_8_adj_2356), .CI(co_mult_10u_9u_0_0_3_adj_2344), 
           .COUT(co_mult_10u_9u_0_0_4_adj_2351), .S0(s_mult_10u_9u_0_0_7_adj_2352), 
           .S1(s_mult_10u_9u_0_0_8_adj_2353)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_0_5_adj_534 (.A0(mult_10u_9u_0_pp_0_9_adj_2362), 
           .A1(mult_10u_9u_0_pp_0_10_adj_2361), .B0(mult_10u_9u_0_pp_1_9_adj_2364), 
           .B1(mult_10u_9u_0_pp_1_10_adj_2363), .CI(co_mult_10u_9u_0_0_4_adj_2351), 
           .COUT(co_mult_10u_9u_0_0_5_adj_2358), .S0(s_mult_10u_9u_0_0_9_adj_2359), 
           .S1(s_mult_10u_9u_0_0_10_adj_2360)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_0_6_adj_535 (.A0(mult_10u_9u_0_pp_0_11_adj_2325), 
           .A1(GND_net), .B0(mult_10u_9u_0_pp_1_11_adj_2369), .B1(mult_10u_9u_0_pp_1_12_adj_2368), 
           .CI(co_mult_10u_9u_0_0_5_adj_2358), .COUT(co_mult_10u_9u_0_0_6_adj_2365), 
           .S0(s_mult_10u_9u_0_0_11_adj_2366), .S1(s_mult_10u_9u_0_0_12_adj_2367)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_0_7_adj_536 (.A0(GND_net), .A1(GND_net), .B0(mult_10u_9u_0_pp_1_13_adj_2328), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_0_6_adj_2365), .COUT(co_mult_10u_9u_0_0_7_adj_2370), 
           .S0(s_mult_10u_9u_0_0_13_adj_2371), .S1(s_mult_10u_9u_0_0_14_adj_2372)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B Cadd_mult_10u_9u_0_0_8_adj_537 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_0_7_adj_2370), .S0(s_mult_10u_9u_0_0_15_adj_2373)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B Cadd_mult_10u_9u_0_1_1_adj_538 (.A0(GND_net), .A1(mult_10u_9u_0_pp_2_6_adj_2376), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_3_6_adj_2322), .CI(GND_net), 
           .COUT(co_mult_10u_9u_0_1_1_adj_2374), .S1(s_mult_10u_9u_0_1_6_adj_2375)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_1_2_adj_539 (.A0(mult_10u_9u_0_pp_2_7_adj_2381), 
           .A1(mult_10u_9u_0_pp_2_8_adj_2380), .B0(mult_10u_9u_0_pp_3_7_adj_2383), 
           .B1(mult_10u_9u_0_pp_3_8_adj_2382), .CI(co_mult_10u_9u_0_1_1_adj_2374), 
           .COUT(co_mult_10u_9u_0_1_2_adj_2377), .S0(s_mult_10u_9u_0_1_7_adj_2378), 
           .S1(s_mult_10u_9u_0_1_8_adj_2379)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_1_3_adj_540 (.A0(mult_10u_9u_0_pp_2_9_adj_2388), 
           .A1(mult_10u_9u_0_pp_2_10_adj_2387), .B0(mult_10u_9u_0_pp_3_9_adj_2390), 
           .B1(mult_10u_9u_0_pp_3_10_adj_2389), .CI(co_mult_10u_9u_0_1_2_adj_2377), 
           .COUT(co_mult_10u_9u_0_1_3_adj_2384), .S0(s_mult_10u_9u_0_1_9_adj_2385), 
           .S1(s_mult_10u_9u_0_1_10_adj_2386)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_1_4_adj_541 (.A0(mult_10u_9u_0_pp_2_11_adj_2395), 
           .A1(mult_10u_9u_0_pp_2_12_adj_2394), .B0(mult_10u_9u_0_pp_3_11_adj_2397), 
           .B1(mult_10u_9u_0_pp_3_12_adj_2396), .CI(co_mult_10u_9u_0_1_3_adj_2384), 
           .COUT(co_mult_10u_9u_0_1_4_adj_2391), .S0(s_mult_10u_9u_0_1_11_adj_2392), 
           .S1(s_mult_10u_9u_0_1_12_adj_2393)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_1_5_adj_542 (.A0(mult_10u_9u_0_pp_2_13_adj_2402), 
           .A1(mult_10u_9u_0_pp_2_14_adj_2401), .B0(mult_10u_9u_0_pp_3_13_adj_2404), 
           .B1(mult_10u_9u_0_pp_3_14_adj_2403), .CI(co_mult_10u_9u_0_1_4_adj_2391), 
           .COUT(co_mult_10u_9u_0_1_5_adj_2398), .S0(s_mult_10u_9u_0_1_13_adj_2399), 
           .S1(s_mult_10u_9u_0_1_14_adj_2400)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_1_6_adj_543 (.A0(mult_10u_9u_0_pp_2_15_adj_2331), 
           .A1(GND_net), .B0(mult_10u_9u_0_pp_3_15_adj_2409), .B1(mult_10u_9u_0_pp_3_16_adj_2408), 
           .CI(co_mult_10u_9u_0_1_5_adj_2398), .COUT(co_mult_10u_9u_0_1_6_adj_2405), 
           .S0(s_mult_10u_9u_0_1_15_adj_2406), .S1(s_mult_10u_9u_0_1_16_adj_2407)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_1_7_adj_544 (.A0(GND_net), .A1(GND_net), .B0(mult_10u_9u_0_pp_3_17_adj_2334), 
           .B1(GND_net), .CI(co_mult_10u_9u_0_1_6_adj_2405), .S0(s_mult_10u_9u_0_1_17_adj_2410), 
           .S1(s_mult_10u_9u_0_1_18_adj_2411)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B Cadd_mult_10u_9u_0_2_1_adj_545 (.A0(GND_net), .A1(s_mult_10u_9u_0_0_4_adj_2339), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_2_4_adj_2323), .CI(GND_net), 
           .COUT(co_mult_10u_9u_0_2_1_adj_2412), .S1(RED_OUT_9__N_613[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_2_adj_546 (.A0(s_mult_10u_9u_0_0_5_adj_2345), 
           .A1(s_mult_10u_9u_0_0_6_adj_2346), .B0(mult_10u_9u_0_pp_2_5_adj_2414), 
           .B1(s_mult_10u_9u_0_1_6_adj_2375), .CI(co_mult_10u_9u_0_2_1_adj_2412), 
           .COUT(co_mult_10u_9u_0_2_2_adj_2413), .S0(RED_OUT_9__N_613[5]), 
           .S1(RED_OUT_9__N_613[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_3_adj_547 (.A0(s_mult_10u_9u_0_0_7_adj_2352), 
           .A1(s_mult_10u_9u_0_0_8_adj_2353), .B0(s_mult_10u_9u_0_1_7_adj_2378), 
           .B1(s_mult_10u_9u_0_1_8_adj_2379), .CI(co_mult_10u_9u_0_2_2_adj_2413), 
           .COUT(co_mult_10u_9u_0_2_3_adj_2415), .S0(RED_OUT_9__N_613[7]), 
           .S1(s_mult_10u_9u_0_2_8_adj_2416)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_4_adj_548 (.A0(s_mult_10u_9u_0_0_9_adj_2359), 
           .A1(s_mult_10u_9u_0_0_10_adj_2360), .B0(s_mult_10u_9u_0_1_9_adj_2385), 
           .B1(s_mult_10u_9u_0_1_10_adj_2386), .CI(co_mult_10u_9u_0_2_3_adj_2415), 
           .COUT(co_mult_10u_9u_0_2_4_adj_2417), .S0(s_mult_10u_9u_0_2_9_adj_2418), 
           .S1(s_mult_10u_9u_0_2_10_adj_2419)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_5_adj_549 (.A0(s_mult_10u_9u_0_0_11_adj_2366), 
           .A1(s_mult_10u_9u_0_0_12_adj_2367), .B0(s_mult_10u_9u_0_1_11_adj_2392), 
           .B1(s_mult_10u_9u_0_1_12_adj_2393), .CI(co_mult_10u_9u_0_2_4_adj_2417), 
           .COUT(co_mult_10u_9u_0_2_5_adj_2420), .S0(s_mult_10u_9u_0_2_11_adj_2421), 
           .S1(s_mult_10u_9u_0_2_12_adj_2422)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_6_adj_550 (.A0(s_mult_10u_9u_0_0_13_adj_2371), 
           .A1(s_mult_10u_9u_0_0_14_adj_2372), .B0(s_mult_10u_9u_0_1_13_adj_2399), 
           .B1(s_mult_10u_9u_0_1_14_adj_2400), .CI(co_mult_10u_9u_0_2_5_adj_2420), 
           .COUT(co_mult_10u_9u_0_2_6_adj_2423), .S0(s_mult_10u_9u_0_2_13_adj_2424), 
           .S1(s_mult_10u_9u_0_2_14_adj_2425)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_7_adj_551 (.A0(s_mult_10u_9u_0_0_15_adj_2373), 
           .A1(GND_net), .B0(s_mult_10u_9u_0_1_15_adj_2406), .B1(s_mult_10u_9u_0_1_16_adj_2407), 
           .CI(co_mult_10u_9u_0_2_6_adj_2423), .COUT(co_mult_10u_9u_0_2_7_adj_2426), 
           .S0(s_mult_10u_9u_0_2_15_adj_2427), .S1(s_mult_10u_9u_0_2_16_adj_2428)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B mult_10u_9u_0_add_2_8_adj_552 (.A0(GND_net), .A1(GND_net), .B0(s_mult_10u_9u_0_1_17_adj_2410), 
           .B1(s_mult_10u_9u_0_1_18_adj_2411), .CI(co_mult_10u_9u_0_2_7_adj_2426), 
           .S0(s_mult_10u_9u_0_2_17_adj_2429), .S1(s_mult_10u_9u_0_2_18_adj_2430)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B Cadd_t_mult_10u_9u_0_3_1_adj_553 (.A0(GND_net), .A1(s_mult_10u_9u_0_2_8_adj_2416), 
           .B0(GND_net), .B1(mult_10u_9u_0_pp_4_8_adj_2140), .CI(GND_net), 
           .COUT(co_t_mult_10u_9u_0_3_1_adj_2431), .S1(RED_OUT_9__N_613[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B t_mult_10u_9u_0_add_3_2_adj_554 (.A0(s_mult_10u_9u_0_2_9_adj_2418), 
           .A1(s_mult_10u_9u_0_2_10_adj_2419), .B0(mult_10u_9u_0_pp_4_9_adj_2432), 
           .B1(mult_10u_9u_0_pp_4_10_adj_2433), .CI(co_t_mult_10u_9u_0_3_1_adj_2431), 
           .COUT(co_t_mult_10u_9u_0_3_2_adj_2434), .S0(RED_OUT_9__N_613[9]), 
           .S1(RED_OUT_9__N_613[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B t_mult_10u_9u_0_add_3_3_adj_555 (.A0(s_mult_10u_9u_0_2_11_adj_2421), 
           .A1(s_mult_10u_9u_0_2_12_adj_2422), .B0(mult_10u_9u_0_pp_4_11_adj_2435), 
           .B1(mult_10u_9u_0_pp_4_12_adj_2436), .CI(co_t_mult_10u_9u_0_3_2_adj_2434), 
           .COUT(co_t_mult_10u_9u_0_3_3_adj_2437), .S0(RED_OUT_9__N_613[11]), 
           .S1(RED_OUT_9__N_613[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B t_mult_10u_9u_0_add_3_4_adj_556 (.A0(s_mult_10u_9u_0_2_13_adj_2424), 
           .A1(s_mult_10u_9u_0_2_14_adj_2425), .B0(mult_10u_9u_0_pp_4_13_adj_2438), 
           .B1(mult_10u_9u_0_pp_4_14_adj_2439), .CI(co_t_mult_10u_9u_0_3_3_adj_2437), 
           .COUT(co_t_mult_10u_9u_0_3_4_adj_2440), .S0(RED_OUT_9__N_613[13]), 
           .S1(RED_OUT_9__N_613[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B t_mult_10u_9u_0_add_3_5_adj_557 (.A0(s_mult_10u_9u_0_2_15_adj_2427), 
           .A1(s_mult_10u_9u_0_2_16_adj_2428), .B0(mult_10u_9u_0_pp_4_15_adj_2441), 
           .B1(mult_10u_9u_0_pp_4_16_adj_2442), .CI(co_t_mult_10u_9u_0_3_4_adj_2440), 
           .COUT(co_t_mult_10u_9u_0_3_5_adj_2443), .S0(RED_OUT_9__N_613[15]), 
           .S1(RED_OUT_9__N_613[16])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    FADD2B t_mult_10u_9u_0_add_3_6_adj_558 (.A0(s_mult_10u_9u_0_2_17_adj_2429), 
           .A1(s_mult_10u_9u_0_2_18_adj_2430), .B0(mult_10u_9u_0_pp_4_17_adj_2444), 
           .B1(GND_net), .CI(co_t_mult_10u_9u_0_3_5_adj_2443), .S0(RED_OUT_9__N_613[17]), 
           .S1(RED_OUT_9__N_613[18])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_0_0_adj_559 (.A0(VRAM_DATA_OUT[0]), .A1(VRAM_DATA_OUT[1]), 
          .A2(VRAM_DATA_OUT[1]), .A3(VRAM_DATA_OUT[2]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mult_10u_9u_0_cin_lr_0_adj_2445), .CO(mco_adj_2446), .P0(RED_OUT_9__N_613[1]), 
          .P1(mult_10u_9u_0_pp_0_2_adj_2337)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_0_1_adj_560 (.A0(VRAM_DATA_OUT[2]), .A1(VRAM_DATA_OUT[3]), 
          .A2(VRAM_DATA_OUT[3]), .A3(VRAM_DATA_OUT[4]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_adj_2446), .CO(mco_1_adj_2447), .P0(mult_10u_9u_0_pp_0_3_adj_2341), 
          .P1(mult_10u_9u_0_pp_0_4_adj_2340)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_0_2_adj_561 (.A0(VRAM_DATA_OUT[4]), .A1(VRAM_DATA_OUT[5]), 
          .A2(VRAM_DATA_OUT[5]), .A3(VRAM_DATA_OUT[6]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_1_adj_2447), .CO(mco_2_adj_2448), .P0(mult_10u_9u_0_pp_0_5_adj_2348), 
          .P1(mult_10u_9u_0_pp_0_6_adj_2347)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_0_3_adj_562 (.A0(VRAM_DATA_OUT[6]), .A1(VRAM_DATA_OUT[7]), 
          .A2(VRAM_DATA_OUT[7]), .A3(VRAM_DATA_OUT[8]), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_2_adj_2448), .CO(mco_3_adj_2449), .P0(mult_10u_9u_0_pp_0_7_adj_2355), 
          .P1(mult_10u_9u_0_pp_0_8_adj_2354)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_0_4_adj_563 (.A0(VRAM_DATA_OUT[8]), .A1(VRAM_DATA_OUT[9]), 
          .A2(VRAM_DATA_OUT[9]), .A3(GND_net), .B0(RED_OUT_9__N_768[1]), 
          .B1(RED_OUT_9__N_768[0]), .B2(RED_OUT_9__N_768[1]), .B3(RED_OUT_9__N_768[0]), 
          .CI(mco_3_adj_2449), .CO(mfco_adj_2326), .P0(mult_10u_9u_0_pp_0_9_adj_2362), 
          .P1(mult_10u_9u_0_pp_0_10_adj_2361)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_2_0_adj_564 (.A0(VRAM_DATA_OUT[0]), .A1(VRAM_DATA_OUT[1]), 
          .A2(VRAM_DATA_OUT[1]), .A3(VRAM_DATA_OUT[2]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mult_10u_9u_0_cin_lr_2_adj_2327), .CO(mco_4_adj_2450), .P0(mult_10u_9u_0_pp_1_3_adj_2343), 
          .P1(mult_10u_9u_0_pp_1_4_adj_2342)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_2_1_adj_565 (.A0(VRAM_DATA_OUT[2]), .A1(VRAM_DATA_OUT[3]), 
          .A2(VRAM_DATA_OUT[3]), .A3(VRAM_DATA_OUT[4]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_4_adj_2450), .CO(mco_5_adj_2451), .P0(mult_10u_9u_0_pp_1_5_adj_2350), 
          .P1(mult_10u_9u_0_pp_1_6_adj_2349)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_2_2_adj_566 (.A0(VRAM_DATA_OUT[4]), .A1(VRAM_DATA_OUT[5]), 
          .A2(VRAM_DATA_OUT[5]), .A3(VRAM_DATA_OUT[6]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_5_adj_2451), .CO(mco_6_adj_2452), .P0(mult_10u_9u_0_pp_1_7_adj_2357), 
          .P1(mult_10u_9u_0_pp_1_8_adj_2356)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_2_3_adj_567 (.A0(VRAM_DATA_OUT[6]), .A1(VRAM_DATA_OUT[7]), 
          .A2(VRAM_DATA_OUT[7]), .A3(VRAM_DATA_OUT[8]), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_6_adj_2452), .CO(mco_7_adj_2453), .P0(mult_10u_9u_0_pp_1_9_adj_2364), 
          .P1(mult_10u_9u_0_pp_1_10_adj_2363)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_2_4_adj_568 (.A0(VRAM_DATA_OUT[8]), .A1(VRAM_DATA_OUT[9]), 
          .A2(VRAM_DATA_OUT[9]), .A3(GND_net), .B0(RED_OUT_9__N_768[3]), 
          .B1(RED_OUT_9__N_768[2]), .B2(RED_OUT_9__N_768[3]), .B3(RED_OUT_9__N_768[2]), 
          .CI(mco_7_adj_2453), .CO(mfco_1_adj_2329), .P0(mult_10u_9u_0_pp_1_11_adj_2369), 
          .P1(mult_10u_9u_0_pp_1_12_adj_2368)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_4_0_adj_569 (.A0(VRAM_DATA_OUT[0]), .A1(VRAM_DATA_OUT[1]), 
          .A2(VRAM_DATA_OUT[1]), .A3(VRAM_DATA_OUT[2]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mult_10u_9u_0_cin_lr_4_adj_2330), .CO(mco_8_adj_2454), .P0(mult_10u_9u_0_pp_2_5_adj_2414), 
          .P1(mult_10u_9u_0_pp_2_6_adj_2376)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_4_1_adj_570 (.A0(VRAM_DATA_OUT[2]), .A1(VRAM_DATA_OUT[3]), 
          .A2(VRAM_DATA_OUT[3]), .A3(VRAM_DATA_OUT[4]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_8_adj_2454), .CO(mco_9_adj_2455), .P0(mult_10u_9u_0_pp_2_7_adj_2381), 
          .P1(mult_10u_9u_0_pp_2_8_adj_2380)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_4_2_adj_571 (.A0(VRAM_DATA_OUT[4]), .A1(VRAM_DATA_OUT[5]), 
          .A2(VRAM_DATA_OUT[5]), .A3(VRAM_DATA_OUT[6]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_9_adj_2455), .CO(mco_10_adj_2456), .P0(mult_10u_9u_0_pp_2_9_adj_2388), 
          .P1(mult_10u_9u_0_pp_2_10_adj_2387)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_4_3_adj_572 (.A0(VRAM_DATA_OUT[6]), .A1(VRAM_DATA_OUT[7]), 
          .A2(VRAM_DATA_OUT[7]), .A3(VRAM_DATA_OUT[8]), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_10_adj_2456), .CO(mco_11_adj_2457), .P0(mult_10u_9u_0_pp_2_11_adj_2395), 
          .P1(mult_10u_9u_0_pp_2_12_adj_2394)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_4_4_adj_573 (.A0(VRAM_DATA_OUT[8]), .A1(VRAM_DATA_OUT[9]), 
          .A2(VRAM_DATA_OUT[9]), .A3(GND_net), .B0(RED_OUT_9__N_768[5]), 
          .B1(RED_OUT_9__N_768[4]), .B2(RED_OUT_9__N_768[5]), .B3(RED_OUT_9__N_768[4]), 
          .CI(mco_11_adj_2457), .CO(mfco_2_adj_2332), .P0(mult_10u_9u_0_pp_2_13_adj_2402), 
          .P1(mult_10u_9u_0_pp_2_14_adj_2401)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_6_0_adj_574 (.A0(VRAM_DATA_OUT[0]), .A1(VRAM_DATA_OUT[1]), 
          .A2(VRAM_DATA_OUT[1]), .A3(VRAM_DATA_OUT[2]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mult_10u_9u_0_cin_lr_6_adj_2333), .CO(mco_12_adj_2458), .P0(mult_10u_9u_0_pp_3_7_adj_2383), 
          .P1(mult_10u_9u_0_pp_3_8_adj_2382)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_6_1_adj_575 (.A0(VRAM_DATA_OUT[2]), .A1(VRAM_DATA_OUT[3]), 
          .A2(VRAM_DATA_OUT[3]), .A3(VRAM_DATA_OUT[4]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_12_adj_2458), .CO(mco_13_adj_2459), .P0(mult_10u_9u_0_pp_3_9_adj_2390), 
          .P1(mult_10u_9u_0_pp_3_10_adj_2389)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_6_2_adj_576 (.A0(VRAM_DATA_OUT[4]), .A1(VRAM_DATA_OUT[5]), 
          .A2(VRAM_DATA_OUT[5]), .A3(VRAM_DATA_OUT[6]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_13_adj_2459), .CO(mco_14_adj_2460), .P0(mult_10u_9u_0_pp_3_11_adj_2397), 
          .P1(mult_10u_9u_0_pp_3_12_adj_2396)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_6_3_adj_577 (.A0(VRAM_DATA_OUT[6]), .A1(VRAM_DATA_OUT[7]), 
          .A2(VRAM_DATA_OUT[7]), .A3(VRAM_DATA_OUT[8]), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_14_adj_2460), .CO(mco_15_adj_2461), .P0(mult_10u_9u_0_pp_3_13_adj_2404), 
          .P1(mult_10u_9u_0_pp_3_14_adj_2403)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    MULT2 mult_10u_9u_0_mult_6_4_adj_578 (.A0(VRAM_DATA_OUT[8]), .A1(VRAM_DATA_OUT[9]), 
          .A2(VRAM_DATA_OUT[9]), .A3(GND_net), .B0(RED_OUT_9__N_768[7]), 
          .B1(RED_OUT_9__N_768[6]), .B2(RED_OUT_9__N_768[7]), .B3(RED_OUT_9__N_768[6]), 
          .CI(mco_15_adj_2461), .CO(mfco_3_adj_2335), .P0(mult_10u_9u_0_pp_3_15_adj_2409), 
          .P1(mult_10u_9u_0_pp_3_16_adj_2408)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    AND2 AND2_t8_adj_579 (.A(VRAM_DATA_OUT[1]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_9_adj_2432)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(180[10:64])
    AND2 AND2_t7_adj_580 (.A(VRAM_DATA_OUT[2]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_10_adj_2433)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(182[10:65])
    AND2 AND2_t6_adj_581 (.A(VRAM_DATA_OUT[3]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_11_adj_2435)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(184[10:65])
    AND2 AND2_t5_adj_582 (.A(VRAM_DATA_OUT[4]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_12_adj_2436)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(186[10:65])
    AND2 AND2_t4_adj_583 (.A(VRAM_DATA_OUT[5]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_13_adj_2438)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(188[10:65])
    AND2 AND2_t3_adj_584 (.A(VRAM_DATA_OUT[6]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_14_adj_2439)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(190[10:65])
    AND2 AND2_t2_adj_585 (.A(VRAM_DATA_OUT[7]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_15_adj_2441)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(192[10:65])
    AND2 AND2_t1_adj_586 (.A(VRAM_DATA_OUT[8]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_16_adj_2442)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(194[10:65])
    AND2 AND2_t0_adj_587 (.A(VRAM_DATA_OUT[9]), .B(RED_OUT_9__N_768[8]), 
         .Z(mult_10u_9u_0_pp_4_17_adj_2444)) /* synthesis syn_instantiated=1 */ ;   // mult_10u_9u.v(196[10:65])
    FADD2B mult_10u_9u_0_cin_lr_add_0_adj_588 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_10u_9u_0_cin_lr_0_adj_2445)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[57:99])
    CCU2D GREEN_OUT_9__I_0_16 (.A0(GREEN_OUT_9__N_650[14]), .B0(GREEN_OUT_9__N_669[14]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[15]), .B1(GREEN_OUT_9__N_669[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14045), .COUT(n14046), .S0(GREEN_OUT[5]), 
          .S1(GREEN_OUT[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_16.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_16.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_16.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_16.INJECT1_1 = "NO";
    FD1P3AX currSprite_999__i7 (.D(n37[7]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[7])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i7.GSR = "ENABLED";
    FD1P3AX currSprite_999__i6 (.D(n37[6]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[6])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i6.GSR = "ENABLED";
    FD1P3AX currSprite_999__i5 (.D(n37[5]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[5])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i5.GSR = "ENABLED";
    FD1P3AX currSprite_999__i4 (.D(n37[4]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[4])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i4.GSR = "ENABLED";
    FD1P3AX currSprite_999__i3 (.D(n37[3]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[3])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i3.GSR = "ENABLED";
    FD1P3AX currSprite_999__i2 (.D(n37[2]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[2])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i2.GSR = "ENABLED";
    FD1P3AX currSprite_999__i1 (.D(n37[1]), .SP(LOGIC_CLOCK_enable_88), 
            .CK(LOGIC_CLOCK), .Q(currSprite[1])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currSprite_999__i1.GSR = "ENABLED";
    FD1P3AX currValue_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i1.GSR = "DISABLED";
    PFUMX i12621 (.BLUT(n16281), .ALUT(n16282), .C0(n17334), .Z(Sprite_readData2_15__N_492[3]));
    FD1P3AX currValue_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i2.GSR = "DISABLED";
    FD1P3AX currValue_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i3.GSR = "DISABLED";
    FD1P3AX currValue_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i4.GSR = "DISABLED";
    FD1P3AX currValue_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i5.GSR = "DISABLED";
    FD1P3AX currValue_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i6.GSR = "DISABLED";
    FD1P3AX currValue_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currValue[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currValue_i0_i7.GSR = "DISABLED";
    FD1P3AX xPre__i1 (.D(n3189), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i1.GSR = "ENABLED";
    FD1P3AX xPre__i2 (.D(n3190), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i2.GSR = "ENABLED";
    FD1P3AX xPre__i3 (.D(n3191), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i3.GSR = "ENABLED";
    FD1P3AX xPre__i4 (.D(n3192), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i4.GSR = "ENABLED";
    FD1P3AX xPre__i5 (.D(n3193), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i5.GSR = "ENABLED";
    FD1P3AX xPre__i6 (.D(n3194), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i6.GSR = "ENABLED";
    FD1P3AX xPre__i7 (.D(n3195), .SP(LOGIC_CLOCK_enable_102), .CK(LOGIC_CLOCK), 
            .Q(xPre[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam xPre__i7.GSR = "ENABLED";
    FD1P3AX VRAM_ADDR__i2 (.D(SpriteRead_yInSprite_7__N_597[6]), .SP(LOGIC_CLOCK_enable_110), 
            .CK(LOGIC_CLOCK), .Q(\VRAM_ADDR[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i2.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i3 (.D(n17439), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i3.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i4 (.D(n949[1]), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i4.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i5 (.D(n949[2]), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i5.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i6 (.D(n949[3]), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i6.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i7 (.D(n949[4]), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i7.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i8 (.D(n949[5]), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i8.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i9 (.D(n949[6]), .SP(LOGIC_CLOCK_enable_110), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam VRAM_ADDR__i9.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i1 (.D(currColor[1]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currColor_lat_i0_i1.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i2 (.D(currColor[2]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currColor_lat_i0_i2.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i3 (.D(currColor[3]), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam currColor_lat_i0_i3.GSR = "DISABLED";
    FD1P3AX data_0___i2 (.D(VRAM_DATA_9__N_848[1]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i2.GSR = "DISABLED";
    FD1P3AX data_0___i3 (.D(VRAM_DATA_9__N_848[2]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i3.GSR = "DISABLED";
    FD1P3AX data_0___i4 (.D(VRAM_DATA_9__N_848[3]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i4.GSR = "DISABLED";
    FD1P3AX data_0___i5 (.D(VRAM_DATA_9__N_848[4]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i5.GSR = "DISABLED";
    FD1P3AX data_0___i6 (.D(VRAM_DATA_9__N_848[5]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i6.GSR = "DISABLED";
    FD1P3AX data_0___i7 (.D(VRAM_DATA_9__N_848[6]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i7.GSR = "DISABLED";
    FD1P3AX data_0___i8 (.D(VRAM_DATA_9__N_848[7]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i8.GSR = "DISABLED";
    FD1P3AX data_0___i9 (.D(VRAM_DATA_9__N_848[8]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i9.GSR = "DISABLED";
    FD1P3AX data_0___i10 (.D(VRAM_DATA_9__N_848[9]), .SP(LOGIC_CLOCK_enable_122), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_0___i10.GSR = "DISABLED";
    FD1P3AX data_1___i2 (.D(VRAM_DATA_19__N_858[1]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i2.GSR = "DISABLED";
    FD1P3AX data_1___i3 (.D(VRAM_DATA_19__N_858[2]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i3.GSR = "DISABLED";
    FD1P3AX data_1___i4 (.D(VRAM_DATA_19__N_858[3]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i4.GSR = "DISABLED";
    FD1P3AX data_1___i5 (.D(VRAM_DATA_19__N_858[4]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i5.GSR = "DISABLED";
    FD1P3AX data_1___i6 (.D(VRAM_DATA_19__N_858[5]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i6.GSR = "DISABLED";
    FD1P3AX data_1___i7 (.D(VRAM_DATA_19__N_858[6]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[16])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i7.GSR = "DISABLED";
    FD1P3AX data_1___i8 (.D(VRAM_DATA_19__N_858[7]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[17])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i8.GSR = "DISABLED";
    FD1P3AX data_1___i9 (.D(VRAM_DATA_19__N_858[8]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[18])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i9.GSR = "DISABLED";
    FD1P3AX data_1___i10 (.D(VRAM_DATA_19__N_858[9]), .SP(LOGIC_CLOCK_enable_131), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[19])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_1___i10.GSR = "DISABLED";
    FD1P3AX data_2___i2 (.D(VRAM_DATA_29__N_868[1]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[21])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i2.GSR = "DISABLED";
    FD1P3AX data_2___i3 (.D(VRAM_DATA_29__N_868[2]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[22])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i3.GSR = "DISABLED";
    FD1P3AX data_2___i4 (.D(VRAM_DATA_29__N_868[3]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[23])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i4.GSR = "DISABLED";
    FD1P3AX data_2___i5 (.D(VRAM_DATA_29__N_868[4]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[24])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i5.GSR = "DISABLED";
    FD1P3AX data_2___i6 (.D(VRAM_DATA_29__N_868[5]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[25])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i6.GSR = "DISABLED";
    FD1P3AX data_2___i7 (.D(VRAM_DATA_29__N_868[6]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[26])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i7.GSR = "DISABLED";
    FD1P3AX data_2___i8 (.D(VRAM_DATA_29__N_868[7]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[27])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i8.GSR = "DISABLED";
    FD1P3AX data_2___i9 (.D(VRAM_DATA_29__N_868[8]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[28])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i9.GSR = "DISABLED";
    FD1P3AX data_2___i10 (.D(VRAM_DATA_29__N_868[9]), .SP(LOGIC_CLOCK_enable_140), 
            .CK(LOGIC_CLOCK), .Q(VRAM_DATA[29])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam data_2___i10.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i2 (.D(currAddress[1]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i2.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i3 (.D(currAddress[2]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i3.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i4 (.D(currAddress[3]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[3]_adj_2 )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i4.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i5 (.D(currAddress[4]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i5.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i6 (.D(currAddress[5]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i6.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i7 (.D(currAddress[6]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i7.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i8 (.D(currAddress[7]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i8.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i9 (.D(currAddress[8]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i9.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i10 (.D(currAddress[9]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i10.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i11 (.D(currAddress[10]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[10]_adj_18 )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i11.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i12 (.D(currAddress[11]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[11]_adj_19 )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i12.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i13 (.D(currAddress[12]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i13.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i14 (.D(currAddress[13]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[13] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i14.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i15 (.D(currAddress[14]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[14] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i15.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i16 (.D(currAddress[15]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[15] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i16.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i17 (.D(currAddress[16]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[16] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i17.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i18 (.D(currAddress[17]), .SP(LOGIC_CLOCK_enable_157), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[17] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam BUS_ADDR_INTERNAL__i18.GSR = "DISABLED";
    FD1P3DX BUS_transferState_i2 (.D(BUS_transferState_3__N_443[2]), .SP(LOGIC_CLOCK_enable_158), 
            .CK(LOGIC_CLOCK), .CD(n17276), .Q(BUS_transferState[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam BUS_transferState_i2.GSR = "DISABLED";
    PFUMX i12624 (.BLUT(n16284), .ALUT(n16285), .C0(n17334), .Z(Sprite_readData2_15__N_492[4]));
    CCU2D sub_47_add_2_3 (.A0(xPre[1]), .B0(currSprite_pos[1]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[2]), .B1(currSprite_pos[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n14110), .COUT(n14111), .S0(SpriteRead_xInSprite[1]), 
          .S1(SpriteRead_xInSprite[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(273[43:57])
    defparam sub_47_add_2_3.INIT0 = 16'h5999;
    defparam sub_47_add_2_3.INIT1 = 16'h5999;
    defparam sub_47_add_2_3.INJECT1_0 = "NO";
    defparam sub_47_add_2_3.INJECT1_1 = "NO";
    LUT4 i3_3_lut_3_lut_4_lut (.A(LOGIC_CLOCK_enable_52), .B(n18260), .C(n17291), 
         .D(n17276), .Z(LOGIC_CLOCK_enable_165)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i3_3_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 BUS_DONE_OUT_I_63_2_lut_rep_278 (.A(BUS_DONE_OUT_N_1051), .B(otherData2_15__N_540), 
         .Z(n17286)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(564[11:65])
    defparam BUS_DONE_OUT_I_63_2_lut_rep_278.init = 16'h2222;
    LUT4 state_4__bdd_4_lut (.A(state[5]), .B(\state[1] ), .C(\state[3] ), 
         .D(\state[0] ), .Z(n18256)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam state_4__bdd_4_lut.init = 16'h8000;
    LUT4 SpriteRead_xValid_I_0_2_lut (.A(SpriteRead_xValid_N_1166), .B(SpriteRead_xValid_N_1167), 
         .Z(SpriteRead_xValid)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[32:151])
    defparam SpriteRead_xValid_I_0_2_lut.init = 16'h8888;
    FD1P3AX xOffset_pre_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i1.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i2.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i3.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i4.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i5.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i6.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_165), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam xOffset_pre_i0_i7.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i1.GSR = "DISABLED";
    CCU2D sub_47_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[0]), .B1(currSprite_pos[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n14110), .S1(SpriteRead_xInSprite[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(273[43:57])
    defparam sub_47_add_2_1.INIT0 = 16'h0000;
    defparam sub_47_add_2_1.INIT1 = 16'h5999;
    defparam sub_47_add_2_1.INJECT1_0 = "NO";
    defparam sub_47_add_2_1.INJECT1_1 = "NO";
    LUT4 inv_47_i8_1_lut (.A(ALPHA_READ[7]), .Z(RED_OUT_9__N_768[7])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i8_1_lut.init = 16'h5555;
    CCU2D add_1839_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14109), 
          .S0(currAddress_17__N_724[17]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[112:132])
    defparam add_1839_cout.INIT0 = 16'h0000;
    defparam add_1839_cout.INIT1 = 16'h0000;
    defparam add_1839_cout.INJECT1_0 = "NO";
    defparam add_1839_cout.INJECT1_1 = "NO";
    CCU2D add_1839_8 (.A0(y[7]), .B0(n4_adj_2464), .C0(n14511), .D0(GND_net), 
          .A1(y[7]), .B1(n4_adj_2464), .C1(GND_net), .D1(GND_net), .CIN(n14108), 
          .COUT(n14109), .S0(currAddress_17__N_724[15]), .S1(currAddress_17__N_724[16]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[112:132])
    defparam add_1839_8.INIT0 = 16'h9696;
    defparam add_1839_8.INIT1 = 16'h9666;
    defparam add_1839_8.INJECT1_0 = "NO";
    defparam add_1839_8.INJECT1_1 = "NO";
    PFUMX i12627 (.BLUT(n16287), .ALUT(n16288), .C0(n17334), .Z(Sprite_readData2_15__N_492[5]));
    CCU2D add_1839_6 (.A0(y[5]), .B0(SpriteRead_yInSprite_7__N_597[5]), 
          .C0(y[4]), .D0(GND_net), .A1(SpriteRead_yInSprite_7__N_597[6]), 
          .B1(n4_adj_2465), .C1(n30[5]), .D1(GND_net), .CIN(n14107), 
          .COUT(n14108), .S0(currAddress_17__N_724[13]), .S1(currAddress_17__N_724[14]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[112:132])
    defparam add_1839_6.INIT0 = 16'h9696;
    defparam add_1839_6.INIT1 = 16'h9696;
    defparam add_1839_6.INJECT1_0 = "NO";
    defparam add_1839_6.INJECT1_1 = "NO";
    LUT4 i12456_3_lut (.A(n16116), .B(n16117), .C(otherData2_15__N_540), 
         .Z(otherData2[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12456_3_lut.init = 16'hcaca;
    FD1P3AX yOffset_pre_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i2.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i3.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i4.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i5.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i6.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_172), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam yOffset_pre_i0_i7.GSR = "DISABLED";
    FD1P3AX latchMode_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(latchMode[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam latchMode_i0_i1.GSR = "DISABLED";
    FD1P3AX latchMode_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(latchMode[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam latchMode_i0_i2.GSR = "DISABLED";
    FD1P3AX latchMode_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(latchMode[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam latchMode_i0_i3.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i2 (.D(n17342), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i2.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i3 (.D(n17339), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i3.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i4 (.D(n17333), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i4.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i5 (.D(n17332), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i5.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i6 (.D(n17331), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i6.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i7 (.D(n17321), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i7.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i8 (.D(n17334), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i8.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i9 (.D(n17337), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i9.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i10 (.D(n17325), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i10.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i11 (.D(\BUS_addr[10] ), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i11.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i12 (.D(\BUS_addr[11] ), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i12.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i13 (.D(n17335), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i13.GSR = "DISABLED";
    FD1P3AX Sprite_writeAddr__i14 (.D(n17338), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeAddr[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeAddr__i14.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i1.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i2.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i3.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i4.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i5.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i6.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i7.GSR = "DISABLED";
    FD1P3AX Sprite_writeData_i0_i8 (.D(BUS_data[8]), .SP(LOGIC_CLOCK_enable_196), 
            .CK(LOGIC_CLOCK), .Q(Sprite_writeData[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam Sprite_writeData_i0_i8.GSR = "DISABLED";
    FD1S3AX xOffset_i1 (.D(xOffset_pre[1]), .CK(offsetLatchClockOrd), .Q(xOffset[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i1.GSR = "DISABLED";
    FD1S3AX xOffset_i2 (.D(xOffset_pre[2]), .CK(offsetLatchClockOrd), .Q(\xOffset[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i2.GSR = "DISABLED";
    FD1S3AX xOffset_i3 (.D(xOffset_pre[3]), .CK(offsetLatchClockOrd), .Q(\xOffset[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i3.GSR = "DISABLED";
    FD1S3AX xOffset_i4 (.D(xOffset_pre[4]), .CK(offsetLatchClockOrd), .Q(xOffset_c[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i4.GSR = "DISABLED";
    FD1S3AX xOffset_i5 (.D(xOffset_pre[5]), .CK(offsetLatchClockOrd), .Q(xOffset_c[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i5.GSR = "DISABLED";
    FD1S3AX xOffset_i6 (.D(xOffset_pre[6]), .CK(offsetLatchClockOrd), .Q(xOffset_c[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i6.GSR = "DISABLED";
    FD1S3AX xOffset_i7 (.D(xOffset_pre[7]), .CK(offsetLatchClockOrd), .Q(xOffset_c[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=172, LSE_RLINE=172 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(288[3] 291[10])
    defparam xOffset_i7.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_589 (.A(\state[0] ), .B(n19), .C(n15681), .D(n21), 
         .Z(reset_N_1062)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_589.init = 16'hcecc;
    LUT4 i1_4_lut_adj_590 (.A(reset), .B(n5_adj_2321), .C(n17448), .D(n17450), 
         .Z(n19)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_590.init = 16'haaa8;
    LUT4 i1_2_lut_adj_591 (.A(reset), .B(n17275), .Z(n21)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_591.init = 16'hbbbb;
    LUT4 inv_47_i6_1_lut (.A(ALPHA_READ[5]), .Z(RED_OUT_9__N_768[5])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i6_1_lut.init = 16'h5555;
    LUT4 i3_4_lut_adj_592 (.A(n17428), .B(n14320), .C(n17306), .D(n15352), 
         .Z(LOGIC_CLOCK_enable_81)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_592.init = 16'h8000;
    LUT4 i3_2_lut_3_lut (.A(BUS_DONE_OUT_N_1051), .B(otherData2_15__N_540), 
         .C(n15457), .Z(n9)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(564[11:65])
    defparam i3_2_lut_3_lut.init = 16'hd0d0;
    LUT4 state_0__bdd_4_lut_13364 (.A(state[4]), .B(state[7]), .C(state[5]), 
         .D(state[6]), .Z(n17056)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A ((C+(D))+!B))) */ ;
    defparam state_0__bdd_4_lut_13364.init = 16'h2004;
    LUT4 inv_47_i4_1_lut (.A(ALPHA_READ[3]), .Z(RED_OUT_9__N_768[3])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i4_1_lut.init = 16'h5555;
    LUT4 i852_3_lut_rep_276_4_lut_4_lut (.A(otherData2_15__N_540), .B(n2539), 
         .C(n17428), .D(BUS_DONE_OUT_N_1051), .Z(n17284)) /* synthesis lut_function=(!(A (B)+!A (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(582[11:65])
    defparam i852_3_lut_rep_276_4_lut_4_lut.init = 16'h2722;
    CCU2D add_1839_4 (.A0(y[2]), .B0(y[3]), .C0(GND_net), .D0(GND_net), 
          .A1(y[3]), .B1(y[4]), .C1(GND_net), .D1(GND_net), .CIN(n14106), 
          .COUT(n14107), .S0(currAddress_17__N_724[11]), .S1(currAddress_17__N_724[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[112:132])
    defparam add_1839_4.INIT0 = 16'h5666;
    defparam add_1839_4.INIT1 = 16'h5666;
    defparam add_1839_4.INJECT1_0 = "NO";
    defparam add_1839_4.INJECT1_1 = "NO";
    LUT4 i12029_2_lut_3_lut_3_lut (.A(otherData2_15__N_540), .B(n2539), 
         .C(BUS_DONE_OUT_N_1051), .Z(n15689)) /* synthesis lut_function=(!(A (B)+!A !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(582[11:65])
    defparam i12029_2_lut_3_lut_3_lut.init = 16'h7272;
    LUT4 i1_3_lut_2_lut_3_lut_2_lut (.A(otherData2_15__N_540), .B(n2539), 
         .Z(n17287)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(582[11:65])
    defparam i1_3_lut_2_lut_3_lut_2_lut.init = 16'h2222;
    PFUMX i12630 (.BLUT(n16290), .ALUT(n16291), .C0(n17334), .Z(Sprite_readData2_15__N_492[6]));
    LUT4 i11_4_lut (.A(n17340), .B(n22_adj_2467), .C(n18), .D(n17313), 
         .Z(n1985)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i11_4_lut.init = 16'h0040;
    LUT4 i10_4_lut (.A(n19_adj_2468), .B(n17335), .C(n15655), .D(n17411), 
         .Z(n22_adj_2467)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i10_4_lut.init = 16'h0200;
    PFUMX i12633 (.BLUT(n16293), .ALUT(n16294), .C0(n17334), .Z(Sprite_readData2_15__N_492[7]));
    CCU2D add_1839_2 (.A0(currAddress_17__N_724[8]), .B0(y[1]), .C0(GND_net), 
          .D0(GND_net), .A1(y[1]), .B1(y[2]), .C1(GND_net), .D1(GND_net), 
          .COUT(n14106), .S1(currAddress_17__N_724[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[112:132])
    defparam add_1839_2.INIT0 = 16'h7000;
    defparam add_1839_2.INIT1 = 16'h5666;
    defparam add_1839_2.INJECT1_0 = "NO";
    defparam add_1839_2.INJECT1_1 = "NO";
    LUT4 i6_4_lut_adj_593 (.A(n17376), .B(n15436), .C(n15693), .D(n46_c), 
         .Z(n18)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i6_4_lut_adj_593.init = 16'h0400;
    LUT4 i7_4_lut_adj_594 (.A(n17338), .B(n17337), .C(n17380), .D(\BUS_addr[10] ), 
         .Z(n19_adj_2468)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i7_4_lut_adj_594.init = 16'h0100;
    PFUMX i13365 (.BLUT(n17180), .ALUT(n17179), .C0(n1345), .Z(BUS_transferState_3__N_443[0]));
    LUT4 i2_3_lut_3_lut_4_lut (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), .B(n2642), 
         .C(n6135), .D(n17276), .Z(LOGIC_CLOCK_enable_79)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[8:62])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h0020;
    PFUMX i13414 (.BLUT(n17480), .ALUT(n17481), .C0(state[4]), .Z(n17349));
    LUT4 i12033_4_lut (.A(n17362), .B(n17341), .C(n17355), .D(n17383), 
         .Z(n15693)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12033_4_lut.init = 16'hfffe;
    PFUMX i12639 (.BLUT(n16298), .ALUT(n16299), .C0(n17342), .Z(n16301));
    CCU2D GREEN_OUT_9__I_0_14 (.A0(GREEN_OUT_9__N_650[12]), .B0(GREEN_OUT_9__N_669[12]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[13]), .B1(GREEN_OUT_9__N_669[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14044), .COUT(n14045), .S0(GREEN_OUT[3]), 
          .S1(GREEN_OUT[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_14.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_14.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_14.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_14.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_12 (.A0(GREEN_OUT_9__N_650[10]), .B0(GREEN_OUT_9__N_669[10]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[11]), .B1(GREEN_OUT_9__N_669[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14043), .COUT(n14044), .S0(GREEN_OUT[1]), 
          .S1(GREEN_OUT[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_12.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_12.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_12.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_12.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_10 (.A0(GREEN_OUT_9__N_650[8]), .B0(GREEN_OUT_9__N_669[8]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[9]), .B1(GREEN_OUT_9__N_669[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14042), .COUT(n14043), .S1(GREEN_OUT[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_10.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_10.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_10.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_10.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_8 (.A0(GREEN_OUT_9__N_650[6]), .B0(GREEN_OUT_9__N_669[6]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[7]), .B1(GREEN_OUT_9__N_669[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14041), .COUT(n14042));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_8.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_8.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_8.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_8.INJECT1_1 = "NO";
    PFUMX i12643 (.BLUT(n16303), .ALUT(n16304), .C0(n17334), .Z(Sprite_readData2_15__N_492[8]));
    CCU2D GREEN_OUT_9__I_0_6 (.A0(GREEN_OUT_9__N_650[4]), .B0(GREEN_OUT_9__N_669[4]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[5]), .B1(GREEN_OUT_9__N_669[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14040), .COUT(n14041));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_6.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_6.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_6.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_6.INJECT1_1 = "NO";
    CCU2D xPre_7__I_0_752_4 (.A0(xPre[2]), .B0(\xOffset[2] ), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[3]), .B1(\xOffset[3] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n14012), .COUT(n14013), .S0(x[2]), .S1(x[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(249[25:39])
    defparam xPre_7__I_0_752_4.INIT0 = 16'h5666;
    defparam xPre_7__I_0_752_4.INIT1 = 16'h5666;
    defparam xPre_7__I_0_752_4.INJECT1_0 = "NO";
    defparam xPre_7__I_0_752_4.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_4 (.A0(GREEN_OUT_9__N_650[2]), .B0(GREEN_OUT_9__N_669[2]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[3]), .B1(GREEN_OUT_9__N_669[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14039), .COUT(n14040));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_4.INIT0 = 16'h5666;
    defparam GREEN_OUT_9__I_0_4.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_4.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_4.INJECT1_1 = "NO";
    CCU2D add_10513_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n18273), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12]_adj_14 ), 
          .D1(n18272), .CIN(n13997), .COUT(n13998));
    defparam add_10513_5.INIT0 = 16'h00ce;
    defparam add_10513_5.INIT1 = 16'h00ce;
    defparam add_10513_5.INJECT1_0 = "NO";
    defparam add_10513_5.INJECT1_1 = "NO";
    CCU2D add_10513_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[9]_adj_9 ), .D0(n18268), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n18269), 
          .CIN(n13996), .COUT(n13997));
    defparam add_10513_3.INIT0 = 16'h00ce;
    defparam add_10513_3.INIT1 = 16'h00ce;
    defparam add_10513_3.INJECT1_0 = "NO";
    defparam add_10513_3.INJECT1_1 = "NO";
    CCU2D GREEN_OUT_9__I_0_2 (.A0(GREEN_OUT_9__N_650[0]), .B0(GREEN_OUT_9__N_669[0]), 
          .C0(GND_net), .D0(GND_net), .A1(GREEN_OUT_9__N_650[1]), .B1(GREEN_OUT_9__N_669[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n14039));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(281[38:104])
    defparam GREEN_OUT_9__I_0_2.INIT0 = 16'h7000;
    defparam GREEN_OUT_9__I_0_2.INIT1 = 16'h5666;
    defparam GREEN_OUT_9__I_0_2.INJECT1_0 = "NO";
    defparam GREEN_OUT_9__I_0_2.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_20 (.A0(RED_OUT_9__N_613[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14038), .S0(RED_OUT[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_20.INIT0 = 16'h5aaa;
    defparam RED_OUT_9__I_0_20.INIT1 = 16'h0000;
    defparam RED_OUT_9__I_0_20.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_20.INJECT1_1 = "NO";
    LUT4 i5_3_lut_rep_265_3_lut_4_lut (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), 
         .B(n2642), .C(n10_adj_2469), .D(n17276), .Z(n17273)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[8:62])
    defparam i5_3_lut_rep_265_3_lut_4_lut.init = 16'h00d0;
    LUT4 i19_3_lut_4_lut (.A(currSprite_conf[0]), .B(SpriteRead_xValid_N_1166), 
         .C(SpriteRead_xValid_N_1167), .D(state[4]), .Z(n15611)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(197[9:24])
    defparam i19_3_lut_4_lut.init = 16'hc0aa;
    PFUMX i12646 (.BLUT(n16306), .ALUT(n16307), .C0(n17334), .Z(Sprite_readData2_15__N_508[0]));
    PFUMX i12649 (.BLUT(n16309), .ALUT(n16310), .C0(n17334), .Z(Sprite_readData2_15__N_508[1]));
    LUT4 i1_4_lut_rep_341_then_4_lut (.A(state[5]), .B(n15508), .C(state[7]), 
         .D(state[6]), .Z(n17481)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_rep_341_then_4_lut.init = 16'hffef;
    PFUMX i12652 (.BLUT(n16312), .ALUT(n16313), .C0(n17334), .Z(Sprite_readData2_15__N_508[2]));
    PFUMX i12655 (.BLUT(n16315), .ALUT(n16316), .C0(n17334), .Z(Sprite_readData2_15__N_508[3]));
    PFUMX i12661 (.BLUT(n16320), .ALUT(n16321), .C0(n17342), .Z(n16323));
    LUT4 i12949_4_lut_4_lut (.A(n17295), .B(n11_adj_2470), .C(n10_adj_2471), 
         .D(n4), .Z(n12)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[131:253])
    defparam i12949_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i12951_4_lut_4_lut (.A(n17297), .B(n15725), .C(n12_adj_2473), 
         .D(n4_c), .Z(n14)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam i12951_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i2_3_lut_4_lut_adj_595 (.A(n17305), .B(n17298), .C(n63), .D(n63_adj_20), 
         .Z(n14320)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_595.init = 16'he000;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n17305), .B(n17298), .C(n15369), 
         .D(n17276), .Z(LOGIC_CLOCK_enable_175)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h00e0;
    PFUMX i12665 (.BLUT(n16325), .ALUT(n16326), .C0(n17334), .Z(Sprite_readData2_15__N_508[4]));
    PFUMX i12668 (.BLUT(n16328), .ALUT(n16329), .C0(n17334), .Z(Sprite_readData2_15__N_508[5]));
    CCU2D add_579_1724_add_1_10518_add_1_14 (.A0(n3855[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(n3855[13]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n14087), .S0(n16[12]), .S1(n16[13]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_14.INIT0 = 16'hfaaa;
    defparam add_579_1724_add_1_10518_add_1_14.INIT1 = 16'hfaaa;
    defparam add_579_1724_add_1_10518_add_1_14.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_14.INJECT1_1 = "NO";
    CCU2D add_579_1724_add_1_10518_add_1_12 (.A0(n3855[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(n3855[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n14086), .COUT(n14087), .S0(n16[10]), 
          .S1(n16[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_12.INIT0 = 16'hfaaa;
    defparam add_579_1724_add_1_10518_add_1_12.INIT1 = 16'hfaaa;
    defparam add_579_1724_add_1_10518_add_1_12.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_12.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_18 (.A0(RED_OUT_9__N_613[16]), .B0(RED_OUT_9__N_632[16]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[17]), .B1(RED_OUT_9__N_632[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14037), .COUT(n14038), .S0(RED_OUT[7]), 
          .S1(RED_OUT[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_18.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_18.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_18.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_18.INJECT1_1 = "NO";
    PFUMX i12671 (.BLUT(n16331), .ALUT(n16332), .C0(n17334), .Z(Sprite_readData2_15__N_508[6]));
    PFUMX i12674 (.BLUT(n16334), .ALUT(n16335), .C0(n17334), .Z(Sprite_readData2_15__N_508[7]));
    PFUMX i12677 (.BLUT(n16337), .ALUT(n16338), .C0(n17334), .Z(Sprite_readData2_15__N_508[8]));
    CCU2D add_579_1724_add_1_10518_add_1_10 (.A0(n3855[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(n3855[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14085), .COUT(n14086), .S0(n16[8]), .S1(n16[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_10.INIT0 = 16'hfaaa;
    defparam add_579_1724_add_1_10518_add_1_10.INIT1 = 16'hfaaa;
    defparam add_579_1724_add_1_10518_add_1_10.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_10.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_16 (.A0(RED_OUT_9__N_613[14]), .B0(RED_OUT_9__N_632[14]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[15]), .B1(RED_OUT_9__N_632[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14036), .COUT(n14037), .S0(RED_OUT[5]), 
          .S1(RED_OUT[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_16.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_16.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_16.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_16.INJECT1_1 = "NO";
    CCU2D add_579_1724_add_1_10518_add_1_8 (.A0(SpriteRead_xInSprite[6]), 
          .B0(n3855[6]), .C0(GND_net), .D0(GND_net), .A1(SpriteRead_xInSprite[7]), 
          .B1(n3855[7]), .C1(GND_net), .D1(GND_net), .CIN(n14084), .COUT(n14085), 
          .S0(n16[6]), .S1(n16[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_8.INIT0 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_8.INIT1 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_8.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_8.INJECT1_1 = "NO";
    LUT4 SRAM_WE_N_1255_I_0_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17385), .Z(lastAddress_31__N_1434)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_2_lut_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_596 (.A(n17310), .B(n17302), .C(n17309), 
         .D(n17273), .Z(n4486)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i1_2_lut_3_lut_4_lut_adj_596.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_597 (.A(n17310), .B(n17302), .C(n17308), 
         .D(n17273), .Z(n4520)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i1_2_lut_3_lut_4_lut_adj_597.init = 16'h2000;
    CCU2D add_10513_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14002), 
          .S0(otherData2_15__N_540));
    defparam add_10513_cout.INIT0 = 16'h0000;
    defparam add_10513_cout.INIT1 = 16'h0000;
    defparam add_10513_cout.INJECT1_0 = "NO";
    defparam add_10513_cout.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_14 (.A0(RED_OUT_9__N_613[12]), .B0(RED_OUT_9__N_632[12]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[13]), .B1(RED_OUT_9__N_632[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14035), .COUT(n14036), .S0(RED_OUT[3]), 
          .S1(RED_OUT[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_14.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_14.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_14.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_14.INJECT1_1 = "NO";
    CCU2D add_579_1724_add_1_10518_add_1_6 (.A0(SpriteRead_xInSprite[4]), 
          .B0(n3855[4]), .C0(GND_net), .D0(GND_net), .A1(SpriteRead_xInSprite[5]), 
          .B1(n3855[5]), .C1(GND_net), .D1(GND_net), .CIN(n14083), .COUT(n14084), 
          .S0(n16[4]), .S1(n16[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_6.INIT0 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_6.INIT1 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_6.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_6.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_12 (.A0(RED_OUT_9__N_613[10]), .B0(RED_OUT_9__N_632[10]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[11]), .B1(RED_OUT_9__N_632[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14034), .COUT(n14035), .S0(RED_OUT[1]), 
          .S1(RED_OUT[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_12.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_12.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_12.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_12.INJECT1_1 = "NO";
    CCU2D add_10513_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8]_adj_8 ), 
          .D1(n18267), .COUT(n13996));
    defparam add_10513_1.INIT0 = 16'hF000;
    defparam add_10513_1.INIT1 = 16'h00ce;
    defparam add_10513_1.INJECT1_0 = "NO";
    defparam add_10513_1.INJECT1_1 = "NO";
    CCU2D add_10513_13 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14001), .COUT(n14002));
    defparam add_10513_13.INIT0 = 16'heeee;
    defparam add_10513_13.INIT1 = 16'heeee;
    defparam add_10513_13.INJECT1_0 = "NO";
    defparam add_10513_13.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_10 (.A0(RED_OUT_9__N_613[8]), .B0(RED_OUT_9__N_632[8]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[9]), .B1(RED_OUT_9__N_632[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14033), .COUT(n14034), .S1(RED_OUT[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_10.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_10.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_10.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_10.INJECT1_1 = "NO";
    CCU2D add_579_1724_add_1_10518_add_1_4 (.A0(SpriteRead_xInSprite[2]), 
          .B0(n3855[2]), .C0(GND_net), .D0(GND_net), .A1(SpriteRead_xInSprite[3]), 
          .B1(n3855[3]), .C1(GND_net), .D1(GND_net), .CIN(n14082), .COUT(n14083), 
          .S0(n16[2]), .S1(n16[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_4.INIT0 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_4.INIT1 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_4.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_4.INJECT1_1 = "NO";
    PFUMX i12680 (.BLUT(n16340), .ALUT(n16341), .C0(n17334), .Z(Sprite_readData2_15__N_524[0]));
    CCU2D add_10513_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[17]_adj_5 ), .D0(n18264), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), .D1(lastAddress_31__N_1310), 
          .CIN(n14000), .COUT(n14001));
    defparam add_10513_11.INIT0 = 16'h00ce;
    defparam add_10513_11.INIT1 = 16'hff20;
    defparam add_10513_11.INJECT1_0 = "NO";
    defparam add_10513_11.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_8 (.A0(RED_OUT_9__N_613[6]), .B0(RED_OUT_9__N_632[6]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[7]), .B1(RED_OUT_9__N_632[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14032), .COUT(n14033));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_8.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_8.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_8.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_8.INJECT1_1 = "NO";
    CCU2D add_579_1724_add_1_10518_add_1_2 (.A0(SpriteRead_xInSprite[0]), 
          .B0(n3855[0]), .C0(GND_net), .D0(GND_net), .A1(SpriteRead_xInSprite[1]), 
          .B1(n3855[1]), .C1(GND_net), .D1(GND_net), .COUT(n14082), 
          .S1(n16[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[38:97])
    defparam add_579_1724_add_1_10518_add_1_2.INIT0 = 16'h7000;
    defparam add_579_1724_add_1_10518_add_1_2.INIT1 = 16'h5666;
    defparam add_579_1724_add_1_10518_add_1_2.INJECT1_0 = "NO";
    defparam add_579_1724_add_1_10518_add_1_2.INJECT1_1 = "NO";
    LUT4 i11912_3_lut_4_lut (.A(state[5]), .B(n17388), .C(state[6]), .D(state[4]), 
         .Z(n15403)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i11912_3_lut_4_lut.init = 16'h7fff;
    CCU2D RED_OUT_9__I_0_6 (.A0(RED_OUT_9__N_613[4]), .B0(RED_OUT_9__N_632[4]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[5]), .B1(RED_OUT_9__N_632[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14031), .COUT(n14032));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_6.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_6.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_6.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_6.INJECT1_1 = "NO";
    CCU2D RED_OUT_9__I_0_4 (.A0(RED_OUT_9__N_613[2]), .B0(RED_OUT_9__N_632[2]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[3]), .B1(RED_OUT_9__N_632[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14030), .COUT(n14031));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_4.INIT0 = 16'h5666;
    defparam RED_OUT_9__I_0_4.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_4.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_4.INJECT1_1 = "NO";
    CCU2D add_10513_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15]_adj_16 ), .D0(n18271), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16]_adj_15 ), 
          .D1(n18277), .CIN(n13999), .COUT(n14000));
    defparam add_10513_9.INIT0 = 16'hff31;
    defparam add_10513_9.INIT1 = 16'hff31;
    defparam add_10513_9.INJECT1_0 = "NO";
    defparam add_10513_9.INJECT1_1 = "NO";
    PFUMX i94 (.BLUT(n60_adj_2005), .ALUT(n14339), .C0(state[7]), .Z(n93));
    CCU2D add_10508_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14236), 
          .S0(n2642));
    defparam add_10508_cout.INIT0 = 16'h0000;
    defparam add_10508_cout.INIT1 = 16'h0000;
    defparam add_10508_cout.INJECT1_0 = "NO";
    defparam add_10508_cout.INJECT1_1 = "NO";
    CCU2D add_10508_11 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14235), .COUT(n14236));
    defparam add_10508_11.INIT0 = 16'heeee;
    defparam add_10508_11.INIT1 = 16'heeee;
    defparam add_10508_11.INJECT1_0 = "NO";
    defparam add_10508_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_598 (.A(n17310), .B(n17302), .C(n17327), 
         .D(n17273), .Z(n4521)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i1_2_lut_3_lut_4_lut_adj_598.init = 16'h2000;
    LUT4 i12021_3_lut_4_lut (.A(\state[1] ), .B(n17386), .C(state[7]), 
         .D(state[6]), .Z(n15681)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i12021_3_lut_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_599 (.A(n17310), .B(n17302), .C(n17313), 
         .D(n17273), .Z(n4485)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i1_2_lut_3_lut_4_lut_adj_599.init = 16'h0200;
    LUT4 inv_47_i2_1_lut (.A(ALPHA_READ[1]), .Z(RED_OUT_9__N_768[1])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i2_1_lut.init = 16'h5555;
    LUT4 i11972_2_lut_3_lut (.A(lastReadRow_2_derived_5), .B(n17396), .C(\state[0] ), 
         .Z(n15629)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i11972_2_lut_3_lut.init = 16'hfefe;
    LUT4 Sprite_writeClk_N_1144_bdd_4_lut (.A(Sprite_writeClk_N_1144), .B(n17306), 
         .C(n17428), .D(n17286), .Z(BUS_transferState_3__N_926[1])) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam Sprite_writeClk_N_1144_bdd_4_lut.init = 16'h8380;
    CCU2D RED_OUT_9__I_0_2 (.A0(RED_OUT_9__N_613[0]), .B0(RED_OUT_9__N_632[0]), 
          .C0(GND_net), .D0(GND_net), .A1(RED_OUT_9__N_613[1]), .B1(RED_OUT_9__N_632[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n14030));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(280[36:100])
    defparam RED_OUT_9__I_0_2.INIT0 = 16'h7000;
    defparam RED_OUT_9__I_0_2.INIT1 = 16'h5666;
    defparam RED_OUT_9__I_0_2.INJECT1_0 = "NO";
    defparam RED_OUT_9__I_0_2.INJECT1_1 = "NO";
    CCU2D add_24_8 (.A0(currSprite_pos[6]), .B0(\currSprite_size[6] ), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[7]), .B1(\currSprite_size[7] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14028), .S0(SpriteRead_xValid_N_1168[6]), 
          .S1(SpriteRead_xValid_N_1168[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[81:103])
    defparam add_24_8.INIT0 = 16'h5666;
    defparam add_24_8.INIT1 = 16'h5666;
    defparam add_24_8.INJECT1_0 = "NO";
    defparam add_24_8.INJECT1_1 = "NO";
    LUT4 mux_881_i2_3_lut (.A(currSprite_pos[1]), .B(n972[1]), .C(n3201), 
         .Z(n3189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i2_3_lut.init = 16'hcaca;
    LUT4 mux_881_i3_3_lut (.A(currSprite_pos[2]), .B(n972[2]), .C(n3201), 
         .Z(n3190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i3_3_lut.init = 16'hcaca;
    CCU2D add_10508_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[17]_adj_5 ), .D0(n18264), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), .D1(lastAddress_31__N_1310), 
          .CIN(n14234), .COUT(n14235));
    defparam add_10508_9.INIT0 = 16'h00ce;
    defparam add_10508_9.INIT1 = 16'hff20;
    defparam add_10508_9.INJECT1_0 = "NO";
    defparam add_10508_9.INJECT1_1 = "NO";
    CCU2D add_10508_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15]_adj_16 ), .D0(n18271), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16]_adj_15 ), 
          .D1(n18277), .CIN(n14233), .COUT(n14234));
    defparam add_10508_7.INIT0 = 16'h00ce;
    defparam add_10508_7.INIT1 = 16'h00ce;
    defparam add_10508_7.INJECT1_0 = "NO";
    defparam add_10508_7.INJECT1_1 = "NO";
    LUT4 mux_881_i4_3_lut (.A(currSprite_pos[3]), .B(n972[3]), .C(n3201), 
         .Z(n3191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i4_3_lut.init = 16'hcaca;
    LUT4 SpriteRead_yInSprite_7__N_597_7__I_0_i13_2_lut_rep_287 (.A(SpriteRead_yInSprite_7__N_597[6]), 
         .B(SpriteRead_yValid_N_1158_c[6]), .Z(n17295)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[131:253])
    defparam SpriteRead_yInSprite_7__N_597_7__I_0_i13_2_lut_rep_287.init = 16'h6666;
    CCU2D add_10508_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13]_adj_7 ), .D0(n18266), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14]_adj_3 ), 
          .D1(n18262), .CIN(n14232), .COUT(n14233));
    defparam add_10508_5.INIT0 = 16'h00ce;
    defparam add_10508_5.INIT1 = 16'h00ce;
    defparam add_10508_5.INJECT1_0 = "NO";
    defparam add_10508_5.INJECT1_1 = "NO";
    LUT4 mux_881_i5_3_lut (.A(currSprite_pos[4]), .B(n972[4]), .C(n3201), 
         .Z(n3192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i5_3_lut.init = 16'hcaca;
    LUT4 SpriteRead_yInSprite_7__N_597_7__I_0_i10_3_lut_3_lut (.A(SpriteRead_yInSprite_7__N_597[6]), 
         .B(SpriteRead_yValid_N_1158_c[6]), .C(SpriteRead_yValid_N_1158_c[5]), 
         .Z(n10_adj_2471)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[131:253])
    defparam SpriteRead_yInSprite_7__N_597_7__I_0_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_881_i6_3_lut (.A(currSprite_pos[5]), .B(n972[5]), .C(n3201), 
         .Z(n3193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i6_3_lut.init = 16'hcaca;
    CCU2D add_10508_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n18273), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12]_adj_14 ), 
          .D1(n18272), .CIN(n14231), .COUT(n14232));
    defparam add_10508_3.INIT0 = 16'h00ce;
    defparam add_10508_3.INIT1 = 16'h00ce;
    defparam add_10508_3.INJECT1_0 = "NO";
    defparam add_10508_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_341_else_4_lut (.A(n17388), .B(state[5]), .C(state[7]), 
         .D(state[6]), .Z(n17480)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_rep_341_else_4_lut.init = 16'hffdf;
    LUT4 i13091_2_lut_3_lut (.A(SpriteRead_yInSprite_7__N_597[6]), .B(SpriteRead_yValid_N_1158_c[6]), 
         .C(n16473), .Z(n15743)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[131:253])
    defparam i13091_2_lut_3_lut.init = 16'hf6f6;
    LUT4 mux_881_i7_3_lut (.A(currSprite_pos[6]), .B(n972[6]), .C(n3201), 
         .Z(n3194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i7_3_lut.init = 16'hcaca;
    LUT4 mux_881_i8_3_lut (.A(currSprite_pos[7]), .B(n972[7]), .C(n3201), 
         .Z(n3195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i8_3_lut.init = 16'hcaca;
    CCU2D add_10508_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), 
          .D1(n18269), .COUT(n14231));
    defparam add_10508_1.INIT0 = 16'hF000;
    defparam add_10508_1.INIT1 = 16'h00ce;
    defparam add_10508_1.INJECT1_0 = "NO";
    defparam add_10508_1.INJECT1_1 = "NO";
    LUT4 inv_155_i2_1_lut (.A(xPre[1]), .Z(n949[1])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i2_1_lut.init = 16'h5555;
    LUT4 inv_155_i3_1_lut (.A(xPre[2]), .Z(n949[2])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i3_1_lut.init = 16'h5555;
    LUT4 inv_155_i4_1_lut (.A(xPre[3]), .Z(n949[3])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i4_1_lut.init = 16'h5555;
    LUT4 SRAM_WE_N_1255_I_0_293_2_lut_3_lut_4_lut (.A(n17458), .B(n17411), 
         .C(\BUS_addr[11] ), .D(n18270), .Z(lastAddress_31__N_1401)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam SRAM_WE_N_1255_I_0_293_2_lut_3_lut_4_lut.init = 16'h0f0d;
    LUT4 xPre_7__I_0_i13_2_lut_rep_288 (.A(xPre[6]), .B(SpriteRead_xValid_N_1168[6]), 
         .Z(n17296)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i13_2_lut_rep_288.init = 16'h6666;
    LUT4 i13063_2_lut_3_lut (.A(BUS_transferState[0]), .B(BUS_transferState[1]), 
         .C(BUS_transferState[2]), .Z(Sprite_writeClk_N_1144)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(597[11:35])
    defparam i13063_2_lut_3_lut.init = 16'h0202;
    CCU2D add_24_6 (.A0(currSprite_pos[4]), .B0(\currSprite_size[4] ), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[5]), .B1(\currSprite_size[5] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14027), .COUT(n14028), .S0(SpriteRead_xValid_N_1168[4]), 
          .S1(SpriteRead_xValid_N_1168[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[81:103])
    defparam add_24_6.INIT0 = 16'h5666;
    defparam add_24_6.INIT1 = 16'h5666;
    defparam add_24_6.INJECT1_0 = "NO";
    defparam add_24_6.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_451 (.A(BUS_transferState[1]), .B(BUS_transferState[0]), 
         .Z(n17459)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(565[8:32])
    defparam i1_2_lut_rep_451.init = 16'heeee;
    CCU2D add_10509_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14219), .S1(n2504));
    defparam add_10509_21.INIT0 = 16'heeee;
    defparam add_10509_21.INIT1 = 16'h0000;
    defparam add_10509_21.INJECT1_0 = "NO";
    defparam add_10509_21.INJECT1_1 = "NO";
    LUT4 inv_155_i5_1_lut (.A(xPre[4]), .Z(n949[4])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i5_1_lut.init = 16'h5555;
    CCU2D add_10509_19 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[18] ), .D0(lastAddress_31__N_1310), .A1(\BUS_currGrantID[0] ), 
          .B1(\BUS_currGrantID[1] ), .C1(GND_net), .D1(GND_net), .CIN(n14218), 
          .COUT(n14219));
    defparam add_10509_19.INIT0 = 16'hff20;
    defparam add_10509_19.INIT1 = 16'heeee;
    defparam add_10509_19.INJECT1_0 = "NO";
    defparam add_10509_19.INJECT1_1 = "NO";
    LUT4 SRAM_WE_N_1255_I_0_267_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17375), .D(n18270), .Z(lastAddress_31__N_1336)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_267_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 xPre_7__I_0_i10_3_lut_3_lut (.A(xPre[6]), .B(SpriteRead_xValid_N_1168[6]), 
         .C(SpriteRead_xValid_N_1168[5]), .Z(n10_adj_2475)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 inv_155_i6_1_lut (.A(xPre[5]), .Z(n949[5])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i6_1_lut.init = 16'h5555;
    LUT4 inv_155_i7_1_lut (.A(xPre[6]), .Z(n949[6])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(410[48:67])
    defparam inv_155_i7_1_lut.init = 16'h5555;
    LUT4 i2_2_lut_rep_420_3_lut (.A(BUS_transferState[1]), .B(BUS_transferState[0]), 
         .C(BUS_transferState[2]), .Z(n17428)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(565[8:32])
    defparam i2_2_lut_rep_420_3_lut.init = 16'hfefe;
    LUT4 mux_656_i2_3_lut (.A(GR_RE_DOUT[1]), .B(RED_OUT[1]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i2_3_lut.init = 16'hcaca;
    LUT4 xPre_7__I_0_i15_2_lut_rep_289 (.A(xPre[7]), .B(SpriteRead_xValid_N_1168[7]), 
         .Z(n17297)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i15_2_lut_rep_289.init = 16'h6666;
    LUT4 BUS_DONE_OUT_N_1050_bdd_4_lut_4_lut_2_lut (.A(BUS_transferState[0]), 
         .B(BUS_transferState[2]), .Z(n17179)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(565[8:32])
    defparam BUS_DONE_OUT_N_1050_bdd_4_lut_4_lut_2_lut.init = 16'h1111;
    LUT4 mux_656_i3_3_lut (.A(GR_RE_DOUT[2]), .B(RED_OUT[2]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i3_3_lut.init = 16'hcaca;
    LUT4 i6672_2_lut_rep_452 (.A(\state[1] ), .B(\state[0] ), .Z(n17460)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6672_2_lut_rep_452.init = 16'heeee;
    LUT4 xPre_7__I_0_i12_3_lut_3_lut (.A(xPre[7]), .B(SpriteRead_xValid_N_1168[7]), 
         .C(n10_adj_2475), .Z(n12_adj_2473)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_656_i4_3_lut (.A(GR_RE_DOUT[3]), .B(RED_OUT[3]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i4_3_lut.init = 16'hcaca;
    LUT4 mux_656_i5_3_lut (.A(GR_RE_DOUT[4]), .B(RED_OUT[4]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i5_3_lut.init = 16'hcaca;
    LUT4 i13096_2_lut_3_lut (.A(xPre[7]), .B(SpriteRead_xValid_N_1168[7]), 
         .C(n16478), .Z(n15728)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam i13096_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_600 (.A(\state[1] ), .B(\state[0] ), .C(\state[3] ), 
         .D(state[2]), .Z(n15453)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_600.init = 16'h0100;
    LUT4 mux_656_i6_3_lut (.A(GR_RE_DOUT[5]), .B(RED_OUT[5]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i6_3_lut.init = 16'hcaca;
    CCU2D add_10509_17 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[16]_adj_15 ), .D0(n18277), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[17]_adj_5 ), 
          .D1(n18264), .CIN(n14217), .COUT(n14218));
    defparam add_10509_17.INIT0 = 16'h00ce;
    defparam add_10509_17.INIT1 = 16'h00ce;
    defparam add_10509_17.INJECT1_0 = "NO";
    defparam add_10509_17.INJECT1_1 = "NO";
    LUT4 mux_656_i7_3_lut (.A(GR_RE_DOUT[6]), .B(RED_OUT[6]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i7_3_lut.init = 16'hcaca;
    LUT4 mux_656_i8_3_lut (.A(GR_RE_DOUT[7]), .B(RED_OUT[7]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i8_3_lut.init = 16'hcaca;
    LUT4 i76_2_lut_rep_283_3_lut (.A(n17373), .B(n17304), .C(n17305), 
         .Z(n17291)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(536[10:32])
    defparam i76_2_lut_rep_283_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_394_3_lut (.A(\state[1] ), .B(\state[0] ), .C(state[2]), 
         .Z(n17402)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_394_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_601 (.A(n17373), .B(n17304), .C(n17306), 
         .D(n17305), .Z(n7)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(536[10:32])
    defparam i1_2_lut_3_lut_4_lut_adj_601.init = 16'h0f0e;
    LUT4 mux_656_i9_3_lut (.A(GR_RE_DOUT[8]), .B(RED_OUT[8]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i9_3_lut.init = 16'hcaca;
    LUT4 i6596_2_lut_rep_453 (.A(\state[3] ), .B(state[2]), .Z(n17461)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6596_2_lut_rep_453.init = 16'heeee;
    LUT4 mux_656_i10_3_lut (.A(GR_RE_DOUT[9]), .B(RED_OUT[9]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i10_3_lut.init = 16'hcaca;
    CCU2D add_10509_15 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[14]_adj_3 ), .D0(n18262), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[15]_adj_16 ), 
          .D1(n18271), .CIN(n14216), .COUT(n14217));
    defparam add_10509_15.INIT0 = 16'h00ce;
    defparam add_10509_15.INIT1 = 16'h00ce;
    defparam add_10509_15.INJECT1_0 = "NO";
    defparam add_10509_15.INJECT1_1 = "NO";
    LUT4 offsetLatchClock_I_0_4_lut (.A(LOGIC_CLOCK), .B(latchForce), .C(n15410), 
         .D(n9_adj_2477), .Z(offsetLatchClockOrd)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(254[25:55])
    defparam offsetLatchClock_I_0_4_lut.init = 16'hfcee;
    LUT4 i1_3_lut_adj_602 (.A(latchMode[1]), .B(frameEndClock), .C(latchMode[0]), 
         .Z(n15410)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut_adj_602.init = 16'h0808;
    LUT4 i12196_3_lut (.A(n3968), .B(n3984), .C(currSprite[4]), .Z(n15858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12196_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_421_3_lut (.A(\state[3] ), .B(state[2]), .C(state[5]), 
         .Z(n17429)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_421_3_lut.init = 16'hfefe;
    LUT4 mux_710_i2_3_lut (.A(GR_RE_DOUT[1]), .B(GREEN_OUT[1]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i2_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_603 (.A(latchMode[1]), .B(latchMode[2]), .C(latchMode[0]), 
         .D(latchMode[3]), .Z(n9_adj_2477)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+((D)+!C)))) */ ;
    defparam i2_4_lut_adj_603.init = 16'h0012;
    LUT4 mux_710_i3_3_lut (.A(GR_RE_DOUT[2]), .B(GREEN_OUT[2]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i3_3_lut.init = 16'hcaca;
    LUT4 mux_710_i4_3_lut (.A(GR_RE_DOUT[3]), .B(GREEN_OUT[3]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i4_3_lut.init = 16'hcaca;
    CCU2D add_10509_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[12]_adj_14 ), .D0(n18272), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[13]_adj_7 ), 
          .D1(n18266), .CIN(n14215), .COUT(n14216));
    defparam add_10509_13.INIT0 = 16'h00ce;
    defparam add_10509_13.INIT1 = 16'h00ce;
    defparam add_10509_13.INJECT1_0 = "NO";
    defparam add_10509_13.INJECT1_1 = "NO";
    LUT4 mux_710_i5_3_lut (.A(GR_RE_DOUT[4]), .B(GREEN_OUT[4]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i5_3_lut.init = 16'hcaca;
    CCU2D add_10509_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[10] ), .D0(n18269), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[11] ), .D1(n18273), 
          .CIN(n14214), .COUT(n14215));
    defparam add_10509_11.INIT0 = 16'hff31;
    defparam add_10509_11.INIT1 = 16'h00ce;
    defparam add_10509_11.INJECT1_0 = "NO";
    defparam add_10509_11.INJECT1_1 = "NO";
    CCU2D add_10509_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[8]_adj_8 ), .D0(n18267), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[9]_adj_9 ), 
          .D1(n18268), .CIN(n14213), .COUT(n14214));
    defparam add_10509_9.INIT0 = 16'h00ce;
    defparam add_10509_9.INIT1 = 16'h00ce;
    defparam add_10509_9.INJECT1_0 = "NO";
    defparam add_10509_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_604 (.A(n17373), .B(n17304), .C(n15369), 
         .D(n17305), .Z(LOGIC_CLOCK_enable_4)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(536[10:32])
    defparam i1_2_lut_3_lut_4_lut_adj_604.init = 16'hf0e0;
    LUT4 i13018_2_lut_rep_378_3_lut_4_lut (.A(\state[3] ), .B(state[2]), 
         .C(state[4]), .D(state[5]), .Z(n17386)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i13018_2_lut_rep_378_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_351_2_lut_3_lut_4_lut (.A(\state[3] ), .B(state[2]), 
         .C(state[5]), .D(state[6]), .Z(n17359)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_351_2_lut_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_10509_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[6]_adj_12 ), .D0(n18276), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[7]_adj_13 ), 
          .D1(n18274), .CIN(n14212), .COUT(n14213));
    defparam add_10509_7.INIT0 = 16'h00ce;
    defparam add_10509_7.INIT1 = 16'h00ce;
    defparam add_10509_7.INJECT1_0 = "NO";
    defparam add_10509_7.INJECT1_1 = "NO";
    CCU2D add_24_4 (.A0(currSprite_pos[2]), .B0(\currSprite_size[2] ), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[3]), .B1(\currSprite_size[3] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14026), .COUT(n14027), .S0(SpriteRead_xValid_N_1168[2]), 
          .S1(SpriteRead_xValid_N_1168[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[81:103])
    defparam add_24_4.INIT0 = 16'h5666;
    defparam add_24_4.INIT1 = 16'h5666;
    defparam add_24_4.INJECT1_0 = "NO";
    defparam add_24_4.INJECT1_1 = "NO";
    CCU2D add_10509_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[4]_adj_10 ), .D0(n18275), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[5]_adj_6 ), 
          .D1(n18265), .CIN(n14211), .COUT(n14212));
    defparam add_10509_5.INIT0 = 16'h00ce;
    defparam add_10509_5.INIT1 = 16'h00ce;
    defparam add_10509_5.INJECT1_0 = "NO";
    defparam add_10509_5.INJECT1_1 = "NO";
    CCU2D add_10509_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[2]_adj_4 ), .D0(n18263), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[3] ), .D1(n17409), 
          .CIN(n14210), .COUT(n14211));
    defparam add_10509_3.INIT0 = 16'h00ce;
    defparam add_10509_3.INIT1 = 16'h00ce;
    defparam add_10509_3.INJECT1_0 = "NO";
    defparam add_10509_3.INJECT1_1 = "NO";
    LUT4 GR_WR_DOUT_16_15__I_0_i4_3_lut (.A(GR_WR_DOUT_16[3]), .B(otherData2[3]), 
         .C(n17314), .Z(otherData[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_460 (.A(\state[3] ), .B(state[2]), .Z(n17468)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam i1_2_lut_rep_460.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_605 (.A(\state[3] ), .B(state[2]), .C(state[5]), 
         .D(state[6]), .Z(n8405)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam i1_2_lut_3_lut_4_lut_adj_605.init = 16'h0008;
    LUT4 i2_3_lut_4_lut_adj_606 (.A(\state[3] ), .B(state[2]), .C(state[5]), 
         .D(state[4]), .Z(n14338)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[3] 452[10])
    defparam i2_3_lut_4_lut_adj_606.init = 16'h8000;
    CCU2D add_10509_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n17385), .B1(n17458), .C1(n17423), .D1(n18259), .COUT(n14210));
    defparam add_10509_1.INIT0 = 16'hF000;
    defparam add_10509_1.INIT1 = 16'h4448;
    defparam add_10509_1.INJECT1_0 = "NO";
    defparam add_10509_1.INJECT1_1 = "NO";
    CCU2D add_24_2 (.A0(currSprite_pos[0]), .B0(n17394), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[1]), .B1(\currSprite_size[1] ), 
          .C1(GND_net), .D1(GND_net), .COUT(n14026), .S1(SpriteRead_xValid_N_1168[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[81:103])
    defparam add_24_2.INIT0 = 16'h7000;
    defparam add_24_2.INIT1 = 16'h5666;
    defparam add_24_2.INJECT1_0 = "NO";
    defparam add_24_2.INJECT1_1 = "NO";
    CCU2D add_158_9 (.A0(xPre[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14073), 
          .S0(n972[7]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_158_9.INIT0 = 16'h5aaa;
    defparam add_158_9.INIT1 = 16'h0000;
    defparam add_158_9.INJECT1_0 = "NO";
    defparam add_158_9.INJECT1_1 = "NO";
    LUT4 mux_710_i6_3_lut (.A(GR_RE_DOUT[5]), .B(GREEN_OUT[5]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i6_3_lut.init = 16'hcaca;
    LUT4 mux_710_i7_3_lut (.A(GR_RE_DOUT[6]), .B(GREEN_OUT[6]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i7_3_lut.init = 16'hcaca;
    LUT4 mux_710_i8_3_lut (.A(GR_RE_DOUT[7]), .B(GREEN_OUT[7]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i8_3_lut.init = 16'hcaca;
    LUT4 mux_710_i9_3_lut (.A(GR_RE_DOUT[8]), .B(GREEN_OUT[8]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i9_3_lut.init = 16'hcaca;
    LUT4 mux_710_i10_3_lut (.A(GR_RE_DOUT[9]), .B(GREEN_OUT[9]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i10_3_lut.init = 16'hcaca;
    LUT4 mux_664_i2_3_lut (.A(GR_RE_DOUT[1]), .B(BLUE_OUT[1]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i2_3_lut.init = 16'hcaca;
    LUT4 mux_664_i3_3_lut (.A(GR_RE_DOUT[2]), .B(BLUE_OUT[2]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i3_3_lut.init = 16'hcaca;
    LUT4 mux_664_i4_3_lut (.A(GR_RE_DOUT[3]), .B(BLUE_OUT[3]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i4_3_lut.init = 16'hcaca;
    LUT4 mux_664_i5_3_lut (.A(GR_RE_DOUT[4]), .B(BLUE_OUT[4]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i5_3_lut.init = 16'hcaca;
    LUT4 mux_664_i6_3_lut (.A(GR_RE_DOUT[5]), .B(BLUE_OUT[5]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i6_3_lut.init = 16'hcaca;
    LUT4 SRAM_WE_N_1255_I_0_300_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17375), .D(n18270), .Z(lastAddress_31__N_1422)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_300_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 mux_664_i7_3_lut (.A(GR_RE_DOUT[6]), .B(BLUE_OUT[6]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i7_3_lut.init = 16'hcaca;
    LUT4 mux_664_i8_3_lut (.A(GR_RE_DOUT[7]), .B(BLUE_OUT[7]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i8_3_lut.init = 16'hcaca;
    LUT4 i6784_4_lut (.A(GR_WR_DOUT_16[8]), .B(n17272), .C(otherData2[8]), 
         .D(n17314), .Z(\MDM_data[8] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(461[18:101])
    defparam i6784_4_lut.init = 16'h3022;
    LUT4 mux_664_i9_3_lut (.A(GR_RE_DOUT[8]), .B(BLUE_OUT[8]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i9_3_lut.init = 16'hcaca;
    LUT4 xPre_7__I_0_i11_2_lut_rep_292 (.A(xPre[5]), .B(SpriteRead_xValid_N_1168[5]), 
         .Z(n17300)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i11_2_lut_rep_292.init = 16'h6666;
    LUT4 mux_664_i10_3_lut (.A(GR_RE_DOUT[9]), .B(BLUE_OUT[9]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i10_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut (.A(n1339), .B(BUS_transferState[2]), .C(n1345), .D(n17454), 
         .Z(LOGIC_CLOCK_enable_158)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B (C (D))))) */ ;
    defparam i22_4_lut.init = 16'h0535;
    LUT4 i12463_3_lut (.A(n16123), .B(n16124), .C(otherData2_15__N_540), 
         .Z(otherData2[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12463_3_lut.init = 16'hcaca;
    LUT4 i12063_2_lut_3_lut_4_lut (.A(xPre[5]), .B(SpriteRead_xValid_N_1168[5]), 
         .C(SpriteRead_xValid_N_1168[6]), .D(xPre[6]), .Z(n15725)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam i12063_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 i12195_3_lut (.A(n3933), .B(n3949), .C(currSprite[4]), .Z(n15857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12195_3_lut.init = 16'hcaca;
    LUT4 GR_WR_DOUT_16_15__I_0_i10_4_lut (.A(GR_WR_DOUT_16[9]), .B(Sprite_readData2[9]), 
         .C(n17314), .D(otherData2_15__N_540), .Z(\otherData[9] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i10_4_lut.init = 16'h0aca;
    LUT4 xPre_7__I_0_i9_2_lut_rep_293 (.A(xPre[4]), .B(SpriteRead_xValid_N_1168[4]), 
         .Z(n17301)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i9_2_lut_rep_293.init = 16'h6666;
    LUT4 GR_WR_DOUT_16_15__I_0_i5_3_lut (.A(GR_WR_DOUT_16[4]), .B(otherData2[4]), 
         .C(n17314), .Z(otherData[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 BUS_transferState_3__I_0_779_i3_4_lut (.A(n1230), .B(BUS_transferState_3__N_930[2]), 
         .C(n1345), .D(n15448), .Z(BUS_transferState_3__N_443[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[4] 608[11])
    defparam BUS_transferState_3__I_0_779_i3_4_lut.init = 16'hcac0;
    LUT4 n2539_bdd_4_lut (.A(otherData2_15__N_540), .B(n17428), .C(n14320), 
         .D(n17306), .Z(n17175)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n2539_bdd_4_lut.init = 16'h0080;
    LUT4 xPre_7__I_0_i8_3_lut_3_lut (.A(xPre[4]), .B(SpriteRead_xValid_N_1168[4]), 
         .C(n6_adj_2478), .Z(n8_c)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_3_lut_4_lut_adj_607 (.A(n17443), .B(n17397), .C(n15508), .D(n17405), 
         .Z(n15510)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i1_3_lut_4_lut_adj_607.init = 16'hfef0;
    LUT4 inv_47_i1_1_lut (.A(ALPHA_READ[0]), .Z(RED_OUT_9__N_768[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i1_1_lut.init = 16'h5555;
    LUT4 i1586_2_lut (.A(y[5]), .B(SpriteRead_yInSprite_7__N_597[5]), .Z(n30[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[48:59])
    defparam i1586_2_lut.init = 16'h6666;
    CCU2D add_158_7 (.A0(xPre[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14072), 
          .COUT(n14073), .S0(n972[5]), .S1(n972[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_158_7.INIT0 = 16'h5aaa;
    defparam add_158_7.INIT1 = 16'h5aaa;
    defparam add_158_7.INJECT1_0 = "NO";
    defparam add_158_7.INJECT1_1 = "NO";
    LUT4 i4_4_lut_rep_295 (.A(n7_c), .B(lastReadRow[2]), .C(n6), .D(n17407), 
         .Z(lastReadRow_2_derived_5)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[11:36])
    defparam i4_4_lut_rep_295.init = 16'hfbfe;
    LUT4 lastReadRow_4__I_0_i10_1_lut_4_lut (.A(n7_c), .B(lastReadRow[2]), 
         .C(n6), .D(n17407), .Z(state_7__N_345)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(295[11:36])
    defparam lastReadRow_4__I_0_i10_1_lut_4_lut.init = 16'h0401;
    LUT4 i13110_3_lut_4_lut (.A(n17404), .B(n17405), .C(\state[0] ), .D(n15_adj_2023), 
         .Z(n14406)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i13110_3_lut_4_lut.init = 16'h0100;
    LUT4 BUS_transferState_0__bdd_3_lut (.A(BUS_transferState[0]), .B(BUS_transferState[2]), 
         .C(BUS_transferState[1]), .Z(n6135)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam BUS_transferState_0__bdd_3_lut.init = 16'h1010;
    LUT4 i4_4_lut (.A(n5113), .B(n14320), .C(n18260), .D(n17286), .Z(n10_adj_2469)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0800;
    LUT4 state_0__bdd_4_lut_13729 (.A(\state[0] ), .B(n15_adj_2023), .C(n17404), 
         .D(n17405), .Z(LOGIC_CLOCK_enable_49)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B (C+(D))))) */ ;
    defparam state_0__bdd_4_lut_13729.init = 16'h3335;
    LUT4 i2_3_lut (.A(n17380), .B(n17374), .C(n17375), .Z(n15539)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(536[10:32])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut_adj_608 (.A(n17373), .B(n17328), .C(n17305), .D(n15539), 
         .Z(n6340)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(536[10:32])
    defparam i3_4_lut_adj_608.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_609 (.A(\state[0] ), .B(n17404), .C(n17397), 
         .D(n17443), .Z(n15512)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i1_2_lut_3_lut_4_lut_adj_609.init = 16'hfffd;
    LUT4 lastAddress_i1_i19_3_lut_4_lut (.A(n17458), .B(n17411), .C(SRAM_WE_N_1254), 
         .D(\lastAddress[18] ), .Z(n46)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam lastAddress_i1_i19_3_lut_4_lut.init = 16'hfd0d;
    LUT4 SRAM_WE_N_1255_I_0_303_2_lut_2_lut_3_lut_4_lut_4_lut (.A(n17458), 
         .B(n17411), .C(n18270), .D(n17384), .Z(lastAddress_31__N_1431)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_303_2_lut_2_lut_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 i6812_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17371), .Z(GR_WR_ADDR[3])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6812_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_1255_I_0_287_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17381), .Z(lastAddress_31__N_1383)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_287_2_lut_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 i1599_4_lut_3_lut_4_lut (.A(y[5]), .B(SpriteRead_yInSprite_7__N_597[5]), 
         .C(y[6]), .D(SpriteRead_yInSprite_7__N_597[6]), .Z(n4_adj_2464)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[48:59])
    defparam i1599_4_lut_3_lut_4_lut.init = 16'hf880;
    LUT4 i2_3_lut_4_lut_adj_610 (.A(y[5]), .B(SpriteRead_yInSprite_7__N_597[5]), 
         .C(y[6]), .D(SpriteRead_yInSprite_7__N_597[6]), .Z(n14511)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[48:59])
    defparam i2_3_lut_4_lut_adj_610.init = 16'h8778;
    LUT4 i1_2_lut_3_lut_adj_611 (.A(y[5]), .B(SpriteRead_yInSprite_7__N_597[5]), 
         .C(y[6]), .Z(n4_adj_2465)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[48:59])
    defparam i1_2_lut_3_lut_adj_611.init = 16'h7878;
    LUT4 BUS_DONE_OUT_N_1050_bdd_3_lut_4_lut_4_lut (.A(n17314), .B(BUS_DONE_OUT_N_1051), 
         .C(n17428), .D(otherData2_15__N_540), .Z(n17180)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A ((C+(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(548[11:65])
    defparam BUS_DONE_OUT_N_1050_bdd_3_lut_4_lut_4_lut.init = 16'h020e;
    LUT4 i6816_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17373), .Z(GR_WR_ADDR[7])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6816_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    CCU2D add_158_5 (.A0(xPre[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14071), 
          .COUT(n14072), .S0(n972[3]), .S1(n972[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_158_5.INIT0 = 16'h5aaa;
    defparam add_158_5.INIT1 = 16'h5aaa;
    defparam add_158_5.INJECT1_0 = "NO";
    defparam add_158_5.INJECT1_1 = "NO";
    LUT4 i6813_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17375), .Z(GR_WR_ADDR[4])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6813_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 i7001_2_lut_rep_277_3_lut_4_lut (.A(n17458), .B(n17411), .C(n18260), 
         .D(n2642), .Z(n17285)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C+!(D))) */ ;
    defparam i7001_2_lut_rep_277_3_lut_4_lut.init = 16'hf0fd;
    LUT4 i6815_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17374), .Z(GR_WR_ADDR[6])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6815_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 i6814_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17380), .Z(GR_WR_ADDR[5])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6814_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_1255_I_0_256_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17355), .D(n18270), .Z(lastAddress_31__N_1325)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_256_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    CCU2D add_158_3 (.A0(xPre[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14070), 
          .COUT(n14071), .S0(n972[1]), .S1(n972[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_158_3.INIT0 = 16'h5aaa;
    defparam add_158_3.INIT1 = 16'h5aaa;
    defparam add_158_3.INJECT1_0 = "NO";
    defparam add_158_3.INJECT1_1 = "NO";
    LUT4 SRAM_WE_N_1255_I_0_265_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17374), .D(n18270), .Z(lastAddress_31__N_1334)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_265_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 i13010_4_lut (.A(state[2]), .B(n69), .C(n20), .D(n93), .Z(state_7__N_336[0])) /* synthesis lut_function=(!(A (B+(D))+!A (B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i13010_4_lut.init = 16'h0023;
    LUT4 i1_4_lut_adj_612 (.A(\state[0] ), .B(state[2]), .C(n17406), .D(n14412), 
         .Z(n69)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_4_lut_adj_612.init = 16'h4505;
    LUT4 GR_WR_DOUT_16_15__I_0_i6_3_lut (.A(GR_WR_DOUT_16[5]), .B(otherData2[5]), 
         .C(n17314), .Z(otherData[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 i6586_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17385), .Z(GR_WR_ADDR[0])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6586_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 i21_4_lut (.A(n17257), .B(\state[0] ), .C(state[7]), .D(n4_adj_2141), 
         .Z(n20)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(87[9:14])
    defparam i21_4_lut.init = 16'hca0a;
    LUT4 SRAM_WE_N_1255_I_0_257_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17383), .D(n18270), .Z(lastAddress_31__N_1326)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_257_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 SRAM_WE_N_1255_I_0_294_2_lut_3_lut_4_lut (.A(n17458), .B(n17411), 
         .C(\BUS_addr[10] ), .D(n18270), .Z(lastAddress_31__N_1404)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam SRAM_WE_N_1255_I_0_294_2_lut_3_lut_4_lut.init = 16'h0f0d;
    LUT4 SRAM_WE_N_1255_I_0_264_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17373), .D(n18270), .Z(lastAddress_31__N_1333)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_264_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 xPre_7__I_0_i6_3_lut_3_lut (.A(xPre[3]), .B(SpriteRead_xValid_N_1168[3]), 
         .C(SpriteRead_xValid_N_1168[2]), .Z(n6_adj_2478)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam xPre_7__I_0_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i2_3_lut_adj_613 (.A(state[7]), .B(\state[1] ), .C(n15), .Z(n14412)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i2_3_lut_adj_613.init = 16'hefef;
    LUT4 SRAM_WE_N_1255_I_0_266_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17380), .D(n18270), .Z(lastAddress_31__N_1335)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_266_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 SRAM_WE_N_1255_I_0_261_2_lut_3_lut_4_lut (.A(n17458), .B(n17411), 
         .C(\BUS_addr[10] ), .D(n18270), .Z(lastAddress_31__N_1330)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam SRAM_WE_N_1255_I_0_261_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i7_4_lut_adj_614 (.A(n13), .B(n11_adj_2480), .C(xPre[1]), .D(xPre[7]), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(367[8:20])
    defparam i7_4_lut_adj_614.init = 16'hfeff;
    LUT4 SRAM_WE_N_1255_I_0_299_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17380), .D(n18270), .Z(lastAddress_31__N_1419)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_299_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 i12052_3_lut_4_lut (.A(xPre[3]), .B(SpriteRead_xValid_N_1168[3]), 
         .C(SpriteRead_xValid_N_1168[2]), .D(xPre[2]), .Z(n15714)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam i12052_3_lut_4_lut.init = 16'h9009;
    LUT4 i5_4_lut (.A(xPre[0]), .B(xPre[2]), .C(xPre[6]), .D(xPre[4]), 
         .Z(n13)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(367[8:20])
    defparam i5_4_lut.init = 16'hfffe;
    CCU2D add_158_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n14070), 
          .S1(n972[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_158_1.INIT0 = 16'hF000;
    defparam add_158_1.INIT1 = 16'h5555;
    defparam add_158_1.INJECT1_0 = "NO";
    defparam add_158_1.INJECT1_1 = "NO";
    LUT4 i3_2_lut (.A(xPre[3]), .B(xPre[5]), .Z(n11_adj_2480)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(367[8:20])
    defparam i3_2_lut.init = 16'heeee;
    CCU2D add_617_19 (.A0(currAddress_17__N_724[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14069), .S0(currAddress[17]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_19.INIT0 = 16'h5aaa;
    defparam add_617_19.INIT1 = 16'h0000;
    defparam add_617_19.INJECT1_0 = "NO";
    defparam add_617_19.INJECT1_1 = "NO";
    LUT4 inv_47_i9_1_lut (.A(ALPHA_READ[8]), .Z(RED_OUT_9__N_768[8])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i9_1_lut.init = 16'h5555;
    LUT4 SRAM_WE_N_1255_I_0_295_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17376), .D(n18270), .Z(lastAddress_31__N_1407)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_295_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 i12449_3_lut (.A(n16109), .B(n16110), .C(otherData2_15__N_540), 
         .Z(otherData2[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12449_3_lut.init = 16'hcaca;
    LUT4 GR_WR_DOUT_16_15__I_0_i7_3_lut (.A(GR_WR_DOUT_16[6]), .B(otherData2[6]), 
         .C(n17314), .Z(otherData[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 i6810_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17384), .Z(GR_WR_ADDR[1])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6810_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_1255_I_0_291_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17379), .Z(lastAddress_31__N_1395)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_291_2_lut_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 SRAM_WE_N_1255_I_0_288_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17362), .D(n18270), .Z(lastAddress_31__N_1386)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_288_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 SRAM_WE_N_1255_I_0_262_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17376), .D(n18270), .Z(lastAddress_31__N_1331)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_262_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 SRAM_WE_N_1255_I_0_289_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17355), .D(n18270), .Z(lastAddress_31__N_1389)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_289_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 SRAM_WE_N_1255_I_0_292_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17377), .D(n18270), .Z(lastAddress_31__N_1398)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_292_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 GR_WR_DOUT_16_15__I_0_i8_3_lut (.A(GR_WR_DOUT_16[7]), .B(otherData2[7]), 
         .C(n17314), .Z(otherData[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 SRAM_WE_N_1255_I_0_259_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17377), .D(n18270), .Z(lastAddress_31__N_1328)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_259_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 SRAM_WE_N_1255_I_0_290_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17383), .D(n18270), .Z(lastAddress_31__N_1392)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_290_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 i6811_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), .C(n2642), 
         .D(n17382), .Z(GR_WR_ADDR[2])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i6811_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_1255_I_0_258_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17379), .Z(lastAddress_31__N_1327)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_258_2_lut_3_lut_4_lut_4_lut.init = 16'hfd55;
    CCU2D add_617_17 (.A0(currAddress_17__N_724[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_724[16]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n14068), .COUT(n14069), .S0(currAddress[15]), 
          .S1(currAddress[16]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_17.INIT0 = 16'h5aaa;
    defparam add_617_17.INIT1 = 16'h5aaa;
    defparam add_617_17.INJECT1_0 = "NO";
    defparam add_617_17.INJECT1_1 = "NO";
    PFUMX i12335 (.BLUT(n15995), .ALUT(n15996), .C0(currSprite[5]), .Z(currSprite_pos[5]));
    LUT4 i1_2_lut_3_lut_4_lut_adj_615 (.A(n17334), .B(n17321), .C(n17273), 
         .D(n17310), .Z(n4310)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(577[24:69])
    defparam i1_2_lut_3_lut_4_lut_adj_615.init = 16'h0020;
    LUT4 i1_2_lut_adj_616 (.A(\state[0] ), .B(n23_adj_1904), .Z(n73)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_2_lut_adj_616.init = 16'heeee;
    PFUMX i12338 (.BLUT(n15998), .ALUT(n15999), .C0(currSprite[5]), .Z(currSprite_pos[4]));
    LUT4 SRAM_WE_N_1255_I_0_302_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17382), .Z(lastAddress_31__N_1428)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_302_2_lut_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 SRAM_WE_N_1255_I_0_270_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17384), .Z(lastAddress_31__N_1339)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_270_2_lut_3_lut_4_lut_4_lut.init = 16'hfd55;
    PFUMX i12341 (.BLUT(n16001), .ALUT(n16002), .C0(currSprite[5]), .Z(currSprite_pos[3]));
    LUT4 i1_2_lut_adj_617 (.A(n1), .B(LOGIC_CLOCK_enable_33), .Z(n7210)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_617.init = 16'h4444;
    LUT4 SRAM_WE_N_1255_I_0_263_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17378), .Z(lastAddress_31__N_1332)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_263_2_lut_3_lut_4_lut_4_lut.init = 16'hfd55;
    LUT4 GR_WR_DOUT_16_15__I_0_i2_3_lut (.A(GR_WR_DOUT_16[1]), .B(otherData2[1]), 
         .C(n17314), .Z(otherData[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 SRAM_WE_N_1255_I_0_260_2_lut_3_lut_4_lut (.A(n17458), .B(n17411), 
         .C(\BUS_addr[11] ), .D(n18270), .Z(lastAddress_31__N_1329)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam SRAM_WE_N_1255_I_0_260_2_lut_3_lut_4_lut.init = 16'hf0d0;
    PFUMX i12344 (.BLUT(n16004), .ALUT(n16005), .C0(currSprite[5]), .Z(currSprite_size[13]));
    LUT4 i3_4_lut_adj_618 (.A(currColor[3]), .B(currColor[1]), .C(currColor[2]), 
         .D(currColor[0]), .Z(n1)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i3_4_lut_adj_618.init = 16'hfffb;
    LUT4 SRAM_WE_N_1255_I_0_255_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17362), .D(n18270), .Z(lastAddress_31__N_1324)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_255_2_lut_3_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 GR_WR_DOUT_16_15__I_0_i3_3_lut (.A(GR_WR_DOUT_16[2]), .B(otherData2[2]), 
         .C(n17314), .Z(otherData[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(474[15:73])
    defparam GR_WR_DOUT_16_15__I_0_i3_3_lut.init = 16'hcaca;
    PFUMX i12347 (.BLUT(n16007), .ALUT(n16008), .C0(currSprite[5]), .Z(currSprite_pos[2]));
    LUT4 SRAM_WE_N_1255_I_0_271_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17385), .Z(lastAddress_31__N_1340)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_1255_I_0_271_2_lut_3_lut_4_lut_4_lut.init = 16'hfd55;
    LUT4 SRAM_WE_N_1255_I_0_298_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n17374), .D(n18270), .Z(lastAddress_31__N_1416)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_298_2_lut_3_lut_4_lut_4_lut.init = 16'h0a08;
    PFUMX i12350 (.BLUT(n16010), .ALUT(n16011), .C0(currSprite[5]), .Z(currSprite_pos[14]));
    LUT4 SRAM_WE_N_1255_I_0_296_2_lut_3_lut_4_lut_4_lut (.A(n17458), .B(n17411), 
         .C(n18270), .D(n17378), .Z(lastAddress_31__N_1410)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;
    defparam SRAM_WE_N_1255_I_0_296_2_lut_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 i10529_2_lut (.A(currColor[1]), .B(currColor[0]), .Z(n3[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10529_2_lut.init = 16'h6666;
    LUT4 n15343_bdd_4_lut (.A(n15635), .B(state[2]), .C(\state[3] ), .D(n16632), 
         .Z(n17262)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C (D))+!B !(C))) */ ;
    defparam n15343_bdd_4_lut.init = 16'hc101;
    PFUMX i12353 (.BLUT(n16013), .ALUT(n16014), .C0(currSprite[5]), .Z(currSprite_pos[1]));
    LUT4 i84_4_lut_4_lut_then_3_lut (.A(\state[0] ), .B(SpriteRead_xValid_N_1167), 
         .C(SpriteRead_xValid_N_1166), .Z(n17484)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i84_4_lut_4_lut_then_3_lut.init = 16'h4040;
    PFUMX i12356 (.BLUT(n16016), .ALUT(n16017), .C0(currSprite[5]), .Z(currSprite_pos[9]));
    LUT4 i84_4_lut_4_lut_else_3_lut (.A(\state[0] ), .B(n17275), .C(\state[1] ), 
         .D(state[7]), .Z(n17483)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(373[10:23])
    defparam i84_4_lut_4_lut_else_3_lut.init = 16'haa08;
    CCU2D add_19_8 (.A0(currSprite_pos[14]), .B0(currSprite_size[14]), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[15]), .B1(currSprite_size[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14023), .S0(SpriteRead_yValid_N_1158_c[6]), 
          .S1(SpriteRead_yValid_N_1158_c[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[132:154])
    defparam add_19_8.INIT0 = 16'h5666;
    defparam add_19_8.INIT1 = 16'h5666;
    defparam add_19_8.INJECT1_0 = "NO";
    defparam add_19_8.INJECT1_1 = "NO";
    PFUMX i12359 (.BLUT(n16019), .ALUT(n16020), .C0(currSprite[5]), .Z(currSprite_pos[7]));
    LUT4 i10628_2_lut (.A(currAddress_17__N_724[8]), .B(y[1]), .Z(currAddress_17__N_724[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i10628_2_lut.init = 16'h6666;
    LUT4 i3_3_lut_4_lut (.A(n1985), .B(n17274), .C(n17314), .D(otherData2_15__N_540), 
         .Z(n14584)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i3_3_lut_4_lut.init = 16'hffbf;
    LUT4 n14447_bdd_4_lut (.A(n14447), .B(\state[0] ), .C(state[4]), .D(state[7]), 
         .Z(n16771)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D)))) */ ;
    defparam n14447_bdd_4_lut.init = 16'hc0c4;
    LUT4 i12426_3_lut (.A(n16086), .B(n16087), .C(otherData2_15__N_540), 
         .Z(otherData2[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12426_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_4_lut_adj_619 (.A(n17276), .B(n17285), .C(n63), 
         .D(n17291), .Z(LOGIC_CLOCK_enable_172)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(458[95:155])
    defparam i2_3_lut_4_lut_4_lut_adj_619.init = 16'h0100;
    PFUMX i12362 (.BLUT(n16022), .ALUT(n16023), .C0(currSprite[5]), .Z(currSprite_size[14]));
    LUT4 i13048_3_lut_3_lut (.A(n17349), .B(n17265), .C(n15_adj_2023), 
         .Z(state_7__N_336[7])) /* synthesis lut_function=(!(A (B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i13048_3_lut_3_lut.init = 16'h7f7f;
    LUT4 state_1__bdd_4_lut_13533 (.A(\state[1] ), .B(n17386), .C(n14338), 
         .D(state[6]), .Z(n17268)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam state_1__bdd_4_lut_13533.init = 16'hf088;
    LUT4 i11978_4_lut (.A(n17460), .B(n70), .C(n17283), .D(currSprite_conf[0]), 
         .Z(n15635)) /* synthesis lut_function=(A+(B (C (D))+!B (C+!(D)))) */ ;
    defparam i11978_4_lut.init = 16'hfabb;
    PFUMX i12365 (.BLUT(n16025), .ALUT(n16026), .C0(currSprite[5]), .Z(currSprite_size[11]));
    LUT4 i2_4_lut_adj_620 (.A(n1_adj_2481), .B(n15442), .C(n2), .D(n17460), 
         .Z(LOGIC_CLOCK_enable_88)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;
    defparam i2_4_lut_adj_620.init = 16'h00c8;
    LUT4 i13066_4_lut (.A(n17359), .B(\state[1] ), .C(n3198), .D(n11), 
         .Z(LOGIC_CLOCK_enable_102)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i13066_4_lut.init = 16'h0100;
    LUT4 i5282_3_lut (.A(n23_adj_1904), .B(n8625), .C(\state[0] ), .Z(n8626)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(87[9:14])
    defparam i5282_3_lut.init = 16'hc5c5;
    LUT4 mux_881_i1_3_lut (.A(currSprite_pos[0]), .B(n972[0]), .C(n3201), 
         .Z(n3188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_881_i1_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_621 (.A(n1), .B(n17275), .C(SpriteRead_yInSprite_7__N_597[6]), 
         .D(SpriteRead_yInSprite_7__N_597[5]), .Z(n8625)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i3_4_lut_adj_621.init = 16'hefff;
    LUT4 i2_4_lut_adj_622 (.A(n17404), .B(state[6]), .C(n17_adj_2482), 
         .D(lastReadRow_2_derived_5), .Z(LOGIC_CLOCK_enable_110)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut_adj_622.init = 16'h0010;
    LUT4 i12662_3_lut (.A(n16322), .B(n16323), .C(otherData2_15__N_540), 
         .Z(otherData2[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12662_3_lut.init = 16'hcaca;
    PFUMX i12368 (.BLUT(n16028), .ALUT(n16029), .C0(currSprite[5]), .Z(currSprite_pos[12]));
    PFUMX i12371 (.BLUT(n16031), .ALUT(n16032), .C0(currSprite[5]), .Z(currSprite_pos[8]));
    CCU2D add_19_6 (.A0(currSprite_pos[12]), .B0(currSprite_size[12]), .C0(GND_net), 
          .D0(GND_net), .A1(currSprite_pos[13]), .B1(currSprite_size[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14022), .COUT(n14023), .S0(\SpriteRead_yValid_N_1158[4] ), 
          .S1(SpriteRead_yValid_N_1158_c[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[132:154])
    defparam add_19_6.INIT0 = 16'h5666;
    defparam add_19_6.INIT1 = 16'h5666;
    defparam add_19_6.INJECT1_0 = "NO";
    defparam add_19_6.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_623 (.A(n17302), .B(n17273), .C(n17312), .D(Sprite_pointers_N_1136), 
         .Z(Sprite_pointers_N_1123)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(499[3] 609[10])
    defparam i4_4_lut_adj_623.init = 16'h8000;
    PFUMX i12374 (.BLUT(n16034), .ALUT(n16035), .C0(currSprite[5]), .Z(currSprite_pos[0]));
    PFUMX i12377 (.BLUT(n16037), .ALUT(n16038), .C0(currSprite[5]), .Z(currSprite_pos[11]));
    LUT4 i3693_3_lut_4_lut (.A(\state[0] ), .B(n17361), .C(n17360), .D(n1193), 
         .Z(n7044)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i3693_3_lut_4_lut.init = 16'h2f20;
    PFUMX i12380 (.BLUT(n16040), .ALUT(n16041), .C0(currSprite[5]), .Z(currSprite_pos[13]));
    LUT4 i12640_3_lut (.A(n16300), .B(n16301), .C(otherData2_15__N_540), 
         .Z(otherData2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12640_3_lut.init = 16'hcaca;
    CCU2D add_617_15 (.A0(currAddress_17__N_724[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_724[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n14067), .COUT(n14068), .S0(currAddress[13]), 
          .S1(currAddress[14]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_15.INIT0 = 16'h5aaa;
    defparam add_617_15.INIT1 = 16'h5aaa;
    defparam add_617_15.INJECT1_0 = "NO";
    defparam add_617_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_624 (.A(n17343), .B(n17342), .C(n17327), 
         .D(n17273), .Z(n4416)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(572[13:43])
    defparam i1_2_lut_3_lut_4_lut_adj_624.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_625 (.A(n17343), .B(n17342), .C(n17313), 
         .D(n17273), .Z(n4380)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(572[13:43])
    defparam i1_2_lut_3_lut_4_lut_adj_625.init = 16'h0200;
    LUT4 i12612_3_lut (.A(n16272), .B(n16273), .C(otherData2_15__N_540), 
         .Z(otherData2[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12612_3_lut.init = 16'hcaca;
    LUT4 i12439_3_lut (.A(n16099), .B(n16100), .C(otherData2_15__N_540), 
         .Z(otherData2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12439_3_lut.init = 16'hcaca;
    PFUMX i12383 (.BLUT(n16043), .ALUT(n16044), .C0(currSprite[5]), .Z(currSprite_pos[15]));
    LUT4 i12593_3_lut (.A(n16253), .B(n16254), .C(otherData2_15__N_540), 
         .Z(otherData2[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12593_3_lut.init = 16'hcaca;
    CCU2D add_617_13 (.A0(currAddress_17__N_724[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_724[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n14066), .COUT(n14067), .S0(currAddress[11]), 
          .S1(currAddress[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_13.INIT0 = 16'h5aaa;
    defparam add_617_13.INIT1 = 16'h5aaa;
    defparam add_617_13.INJECT1_0 = "NO";
    defparam add_617_13.INJECT1_1 = "NO";
    PFUMX i12386 (.BLUT(n16046), .ALUT(n16047), .C0(currSprite[5]), .Z(currSprite_pos[10]));
    PFUMX i12389 (.BLUT(n16049), .ALUT(n16050), .C0(currSprite[5]), .Z(currSprite_size[10]));
    LUT4 i2_3_lut_4_lut_4_lut_adj_626 (.A(n17276), .B(n15457), .C(n17306), 
         .D(n17291), .Z(LOGIC_CLOCK_enable_196)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(458[95:155])
    defparam i2_3_lut_4_lut_4_lut_adj_626.init = 16'h4000;
    LUT4 i13095_4_lut (.A(n17296), .B(n17300), .C(n17301), .D(n15714), 
         .Z(n16478)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(269[80:150])
    defparam i13095_4_lut.init = 16'hefee;
    LUT4 i12398_3_lut_rep_386 (.A(n16058), .B(n16059), .C(currSprite[5]), 
         .Z(n17394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12398_3_lut_rep_386.init = 16'hcaca;
    LUT4 i10626_2_lut_4_lut (.A(n16058), .B(n16059), .C(currSprite[5]), 
         .D(currSprite_pos[0]), .Z(SpriteRead_xValid_N_1168[0])) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam i10626_2_lut_4_lut.init = 16'h35ca;
    LUT4 i2_4_lut_adj_627 (.A(n15510), .B(n6157), .C(n15512), .D(VRAM_WC), 
         .Z(n14656)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C)))) */ ;
    defparam i2_4_lut_adj_627.init = 16'h7f5f;
    LUT4 i1_4_lut_adj_628 (.A(n15476), .B(n17406), .C(\state[1] ), .D(n55), 
         .Z(n6157)) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_628.init = 16'h8c88;
    LUT4 i2_4_lut_adj_629 (.A(state[7]), .B(state[4]), .C(state[2]), .D(n16632), 
         .Z(n15476)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i2_4_lut_adj_629.init = 16'h0008;
    LUT4 i71_4_lut (.A(state[7]), .B(\state[0] ), .C(state[4]), .D(state[2]), 
         .Z(n55)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i71_4_lut.init = 16'h2134;
    PFUMX i12392 (.BLUT(n16052), .ALUT(n16053), .C0(currSprite[5]), .Z(currSprite_conf[0]));
    LUT4 i1_rep_140_2_lut (.A(\state[0] ), .B(\state[1] ), .Z(n16632)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_rep_140_2_lut.init = 16'h8888;
    LUT4 i6986_2_lut_rep_286_4_lut (.A(\state[3] ), .B(n17446), .C(state[4]), 
         .D(lastReadRow_2_derived_5), .Z(n17294)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i6986_2_lut_rep_286_4_lut.init = 16'hfffb;
    LUT4 i2_4_lut_adj_630 (.A(n17357), .B(SpriteRead_xValid), .C(\state[1] ), 
         .D(\state[0] ), .Z(LOGIC_CLOCK_enable_18)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i2_4_lut_adj_630.init = 16'h0a08;
    LUT4 SpriteRead_yInSprite_7__N_597_7__I_0_i11_2_lut (.A(SpriteRead_yInSprite_7__N_597[5]), 
         .B(SpriteRead_yValid_N_1158_c[5]), .Z(n11_adj_2470)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[131:253])
    defparam SpriteRead_yInSprite_7__N_597_7__I_0_i11_2_lut.init = 16'h9999;
    LUT4 i13090_4_lut (.A(n11_adj_2470), .B(n17299), .C(n17307), .D(n15549), 
         .Z(n16473)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(268[131:253])
    defparam i13090_4_lut.init = 16'h5557;
    LUT4 i1_3_lut_adj_631 (.A(\state[0] ), .B(n17357), .C(\state[1] ), 
         .Z(LOGIC_CLOCK_enable_19)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_adj_631.init = 16'h4848;
    CCU2D add_617_11 (.A0(currAddress_17__N_724[9]), .B0(currAddress_17__N_742[9]), 
          .C0(GND_net), .D0(GND_net), .A1(currAddress_17__N_724[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14065), .COUT(n14066), 
          .S0(currAddress[9]), .S1(currAddress[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_11.INIT0 = 16'h5666;
    defparam add_617_11.INIT1 = 16'h5aaa;
    defparam add_617_11.INJECT1_0 = "NO";
    defparam add_617_11.INJECT1_1 = "NO";
    CCU2D add_617_9 (.A0(currAddress_17__N_742[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_724[8]), .B1(currAddress_17__N_742[8]), 
          .C1(GND_net), .D1(GND_net), .CIN(n14064), .COUT(n14065), .S0(currAddress[7]), 
          .S1(currAddress[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(251[47:168])
    defparam add_617_9.INIT0 = 16'hfaaa;
    defparam add_617_9.INIT1 = 16'h5666;
    defparam add_617_9.INJECT1_0 = "NO";
    defparam add_617_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_632 (.A(currColor_lat[0]), .B(n15528), .C(state[4]), 
         .D(currColor_lat[1]), .Z(LOGIC_CLOCK_enable_122)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+!(D))))) */ ;
    defparam i1_4_lut_adj_632.init = 16'h3031;
    LUT4 mux_656_i1_3_lut (.A(GR_RE_DOUT[0]), .B(RED_OUT[0]), .C(state[4]), 
         .Z(VRAM_DATA_9__N_848[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_656_i1_3_lut.init = 16'hcaca;
    PFUMX i12395 (.BLUT(n16055), .ALUT(n16056), .C0(currSprite[5]), .Z(currSprite_size[15]));
    PFUMX i12401 (.BLUT(n16061), .ALUT(n16062), .C0(currSprite[5]), .Z(\currSprite_size[1] ));
    LUT4 i3_4_lut_adj_633 (.A(state[4]), .B(n6_adj_2004), .C(lastReadRow_2_derived_5), 
         .D(state[7]), .Z(n15528)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_633.init = 16'hfdfe;
    LUT4 i1_4_lut_adj_634 (.A(currColor_lat[0]), .B(n15528), .C(state[4]), 
         .D(currColor_lat[1]), .Z(LOGIC_CLOCK_enable_131)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i1_4_lut_adj_634.init = 16'h3032;
    LUT4 mux_710_i1_3_lut (.A(GR_RE_DOUT[0]), .B(GREEN_OUT[0]), .C(state[4]), 
         .Z(VRAM_DATA_19__N_858[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_710_i1_3_lut.init = 16'hcaca;
    LUT4 mux_664_i1_3_lut (.A(GR_RE_DOUT[0]), .B(BLUE_OUT[0]), .C(state[4]), 
         .Z(VRAM_DATA_29__N_868[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_664_i1_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_635 (.A(state[2]), .B(n17294), .C(n16632), .D(state[7]), 
         .Z(LOGIC_CLOCK_enable_157)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_635.init = 16'h0010;
    LUT4 i4_4_lut_adj_636 (.A(n7_adj_1886), .B(SpriteRead_yInSprite_7__N_597[6]), 
         .C(n17386), .D(SpriteRead_yInSprite_7__N_597[5]), .Z(n1_adj_2481)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut_adj_636.init = 16'h8000;
    LUT4 i12396_3_lut (.A(n4032), .B(n4048), .C(currSprite[4]), .Z(n16058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12396_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_352_3_lut_4_lut (.A(n17450), .B(n17449), .C(n17443), 
         .D(n17448), .Z(n17360)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i1_2_lut_rep_352_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12397_3_lut (.A(n4067), .B(n4083), .C(currSprite[4]), .Z(n16059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12397_3_lut.init = 16'hcaca;
    LUT4 inv_47_i3_1_lut (.A(ALPHA_READ[2]), .Z(RED_OUT_9__N_768[2])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i3_1_lut.init = 16'h5555;
    LUT4 inv_47_i5_1_lut (.A(ALPHA_READ[4]), .Z(RED_OUT_9__N_768[4])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i5_1_lut.init = 16'h5555;
    LUT4 i10625_2_lut (.A(currSprite_pos[8]), .B(currSprite_size[8]), .Z(\SpriteRead_yValid_N_1158[0] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i10625_2_lut.init = 16'h6666;
    LUT4 inv_47_i7_1_lut (.A(ALPHA_READ[6]), .Z(RED_OUT_9__N_768[6])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(282[58:77])
    defparam inv_47_i7_1_lut.init = 16'h5555;
    LUT4 i5_4_lut_adj_637 (.A(n23_adj_1904), .B(state[7]), .C(n15629), 
         .D(n10025), .Z(LOGIC_CLOCK_enable_27)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i5_4_lut_adj_637.init = 16'h0008;
    PFUMX i12404 (.BLUT(n16064), .ALUT(n16065), .C0(currSprite[5]), .Z(\currSprite_size[2] ));
    LUT4 i6687_2_lut (.A(state[2]), .B(\state[1] ), .Z(n10025)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6687_2_lut.init = 16'heeee;
    LUT4 i2075_2_lut_rep_310_3_lut_4_lut (.A(\state[1] ), .B(n17450), .C(\state[0] ), 
         .D(n17405), .Z(n17318)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(319[10:23])
    defparam i2075_2_lut_rep_310_3_lut_4_lut.init = 16'h0010;
    LUT4 n10344_bdd_4_lut_4_lut (.A(n17342), .B(n6340), .C(n17343), .D(n17285), 
         .Z(n15369)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam n10344_bdd_4_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n17342), .B(n17310), .C(n6250), 
         .D(n17343), .Z(LOGIC_CLOCK_enable_54)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0080;
    PFUMX i12407 (.BLUT(n16067), .ALUT(n16068), .C0(currSprite[5]), .Z(\currSprite_size[3] ));
    PFUMX i12410 (.BLUT(n16070), .ALUT(n16071), .C0(currSprite[5]), .Z(\currSprite_size[4] ));
    PFUMX i12413 (.BLUT(n16073), .ALUT(n16074), .C0(currSprite[5]), .Z(\currSprite_size[5] ));
    LUT4 i12_4_lut (.A(n1339), .B(BUS_transferState[2]), .C(n1345), .D(n16805), 
         .Z(LOGIC_CLOCK_enable_48)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B (C (D))))) */ ;
    defparam i12_4_lut.init = 16'h0535;
    LUT4 i1_4_lut_adj_638 (.A(LOGIC_CLOCK_enable_52), .B(n15448), .C(n14320), 
         .D(n17287), .Z(n1345)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_638.init = 16'heaaa;
    PFUMX i12416 (.BLUT(n16076), .ALUT(n16077), .C0(currSprite[5]), .Z(\currSprite_size[6] ));
    LUT4 i1_4_lut_adj_639 (.A(n17284), .B(n14320), .C(BUS_transferState_3__N_930[2]), 
         .D(n17306), .Z(n1339)) /* synthesis lut_function=(A ((C (D))+!B)+!A ((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_639.init = 16'hf377;
    PFUMX i12419 (.BLUT(n16079), .ALUT(n16080), .C0(currSprite[5]), .Z(\currSprite_size[7] ));
    LUT4 equal_695_i13_2_lut_rep_353_3_lut_4_lut (.A(n17448), .B(n17447), 
         .C(n17450), .D(\state[1] ), .Z(n17361)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[7:20])
    defparam equal_695_i13_2_lut_rep_353_3_lut_4_lut.init = 16'hfffe;
    PFUMX i12429 (.BLUT(n16089), .ALUT(n16090), .C0(currSprite[5]), .Z(currSprite_size[8]));
    LUT4 i1_4_lut_adj_640 (.A(n17271), .B(LOGIC_CLOCK_enable_13), .C(n17360), 
         .D(n17318), .Z(LOGIC_CLOCK_enable_29)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_640.init = 16'h8ccc;
    LUT4 i6904_3_lut (.A(SpriteRead_yInSprite_7__N_597[6]), .B(n7044), .C(SpriteRead_yInSprite_7__N_597[5]), 
         .Z(n2194[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i6904_3_lut.init = 16'h4848;
    PFUMX i12432 (.BLUT(n16092), .ALUT(n16093), .C0(currSprite[5]), .Z(currSprite_size[9]));
    LUT4 i13007_4_lut_rep_267 (.A(MDM_done), .B(n15571), .C(n8_adj_21), 
         .D(WRITE_DONE), .Z(n17275)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i13007_4_lut_rep_267.init = 16'h0001;
    LUT4 state_7__I_0_764_i15_2_lut_3_lut_4_lut (.A(n17448), .B(n17447), 
         .C(n17449), .D(n17450), .Z(n15_adj_2082)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[7:20])
    defparam state_7__I_0_764_i15_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_641 (.A(n70), .B(state[5]), .C(n17461), .D(n15611), 
         .Z(n2)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_4_lut_adj_641.init = 16'h0002;
    PFUMX i12442 (.BLUT(n16102), .ALUT(n16103), .C0(currSprite[5]), .Z(currSprite_size[12]));
    LUT4 i7085_2_lut_3_lut_4_lut (.A(\state[3] ), .B(n17446), .C(state[4]), 
         .D(\state[1] ), .Z(n10444)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i7085_2_lut_3_lut_4_lut.init = 16'hf0b0;
    LUT4 i6882_4_lut_4_lut (.A(n17342), .B(n17343), .C(yOffset_c[4]), 
         .D(xOffset_c[4]), .Z(n2872[4])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i6882_4_lut_4_lut.init = 16'h5140;
    LUT4 i1_2_lut_3_lut_4_lut_adj_642 (.A(\state[0] ), .B(n17451), .C(state[2]), 
         .D(\state[3] ), .Z(n70_adj_2484)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_2_lut_3_lut_4_lut_adj_642.init = 16'h8f0f;
    LUT4 i1_2_lut_rep_362_3_lut (.A(\state[0] ), .B(n17451), .C(\state[3] ), 
         .Z(n17370)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i1_2_lut_rep_362_3_lut.init = 16'h8080;
    LUT4 i6883_4_lut_4_lut (.A(n17342), .B(n17343), .C(yOffset_c[5]), 
         .D(xOffset_c[5]), .Z(n2872[5])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i6883_4_lut_4_lut.init = 16'h5140;
    LUT4 i6884_4_lut_4_lut (.A(n17342), .B(n17343), .C(yOffset_c[6]), 
         .D(xOffset_c[6]), .Z(n2872[6])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i6884_4_lut_4_lut.init = 16'h5140;
    LUT4 i1968_4_lut (.A(n5146), .B(n5113), .C(LOGIC_CLOCK_enable_52), 
         .D(n14320), .Z(LOGIC_CLOCK_enable_32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[4] 608[11])
    defparam i1968_4_lut.init = 16'hcacf;
    LUT4 i6885_4_lut_4_lut (.A(n17342), .B(n17343), .C(yOffset_c[7]), 
         .D(xOffset_c[7]), .Z(n2872[7])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 110[10])
    defparam i6885_4_lut_4_lut.init = 16'h5140;
    LUT4 i1961_4_lut (.A(n15689), .B(n6135), .C(n17306), .D(n5113), 
         .Z(n5146)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(511[4] 608[11])
    defparam i1961_4_lut.init = 16'hcac0;
    LUT4 i2_4_lut_adj_643 (.A(n6187), .B(n17446), .C(n15453), .D(state[4]), 
         .Z(n62_adj_1885)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i2_4_lut_adj_643.init = 16'hc088;
    LUT4 i66_4_lut (.A(state[4]), .B(\state[0] ), .C(n70_adj_2484), .D(n10461), 
         .Z(n58)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(87[9:14])
    defparam i66_4_lut.init = 16'ha0b3;
    LUT4 i10527_1_lut (.A(currColor[0]), .Z(n3[0])) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i10527_1_lut.init = 16'h5555;
    LUT4 i7100_3_lut (.A(\state[1] ), .B(state[2]), .C(n17396), .Z(n10461)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i7100_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_644 (.A(LOGIC_CLOCK_enable_52), .B(n6340), .C(n17428), 
         .D(n10346), .Z(n15457)) /* synthesis lut_function=(!(A+(B (C)+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_644.init = 16'h0504;
    LUT4 i1_2_lut_rep_321_3_lut_4_lut (.A(\BUS_ADDR_INTERNAL[1] ), .B(n17456), 
         .C(n17385), .D(n18259), .Z(n17329)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam i1_2_lut_rep_321_3_lut_4_lut.init = 16'hfff8;
    LUT4 otherData_15__N_438_I_0_2_lut_rep_298_4_lut (.A(n17458), .B(n17411), 
         .C(n17344), .D(BUS_DONE_OUT_N_1051), .Z(n17306)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (D))) */ ;
    defparam otherData_15__N_438_I_0_2_lut_rep_298_4_lut.init = 16'h00d5;
    PFUMX i13408 (.BLUT(n17471), .ALUT(n17472), .C0(\BUS_ADDR_INTERNAL[3]_adj_2 ), 
          .Z(n17328));
    LUT4 i6626_2_lut_rep_333_3_lut_4_lut (.A(\BUS_ADDR_INTERNAL[1] ), .B(n17456), 
         .C(n17385), .D(n18259), .Z(n17341)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam i6626_2_lut_rep_333_3_lut_4_lut.init = 16'hf080;
    LUT4 i95_4_lut (.A(\state[0] ), .B(n17370), .C(state[2]), .D(n10444), 
         .Z(n59)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(313[4] 450[11])
    defparam i95_4_lut.init = 16'hc0c5;
    LUT4 i1_2_lut_rep_320_3_lut_4_lut_else_4_lut (.A(n17382), .B(\BUS_ADDR_INTERNAL[3] ), 
         .C(\BUS_currGrantID[1] ), .D(\BUS_currGrantID[0] ), .Z(n17471)) /* synthesis lut_function=(A+!(((D)+!C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(462[18:73])
    defparam i1_2_lut_rep_320_3_lut_4_lut_else_4_lut.init = 16'haaea;
    PFUMX mux_707_i1 (.BLUT(n898[0]), .ALUT(n2191[0]), .C0(n17360), .Z(n2194[0]));
    PFUMX i13132 (.BLUT(n16772), .ALUT(n16771), .C0(\state[1] ), .Z(n16773));
    PFUMX i28 (.BLUT(n15420), .ALUT(n14_adj_2075), .C0(state[7]), .Z(n17_adj_2482));
    SpriteRam SRam (.\Sprite_writeAddr[9] (Sprite_writeAddr[9]), .\Sprite_writeAddr[8] (Sprite_writeAddr[8]), 
            .\Sprite_writeAddr[7] (Sprite_writeAddr[7]), .\Sprite_writeAddr[6] (Sprite_writeAddr[6]), 
            .\Sprite_writeAddr[5] (Sprite_writeAddr[5]), .\Sprite_writeAddr[4] (Sprite_writeAddr[4]), 
            .\Sprite_writeAddr[3] (Sprite_writeAddr[3]), .\Sprite_writeAddr[2] (Sprite_writeAddr[2]), 
            .\Sprite_writeAddr[1] (Sprite_writeAddr[1]), .\Sprite_writeAddr[0] (Sprite_writeAddr[0]), 
            .\Sprite_readAddr[9] (Sprite_readAddr[9]), .\Sprite_readAddr[8] (Sprite_readAddr[8]), 
            .\Sprite_readAddr[7] (Sprite_readAddr[7]), .\Sprite_readAddr[6] (Sprite_readAddr[6]), 
            .\Sprite_readAddr[5] (Sprite_readAddr[5]), .\Sprite_readAddr[4] (Sprite_readAddr[4]), 
            .\Sprite_readAddr[3] (Sprite_readAddr[3]), .\Sprite_readAddr[2] (Sprite_readAddr[2]), 
            .\Sprite_readAddr[1] (Sprite_readAddr[1]), .\Sprite_readAddr[0] (Sprite_readAddr[0]), 
            .Sprite_writeData({Sprite_writeData}), .VCC_net(VCC_net), .Sprite_readClk(Sprite_readClk), 
            .GND_net(GND_net), .Sprite_writeClk(Sprite_writeClk), .\Sprite_readAddr[11] (Sprite_readAddr[11]), 
            .\Sprite_readAddr[12] (Sprite_readAddr[12]), .\Sprite_readAddr[13] (Sprite_readAddr[13]), 
            .\Sprite_writeAddr[11] (Sprite_writeAddr[11]), .\Sprite_writeAddr[10] (Sprite_writeAddr[10]), 
            .\Sprite_writeAddr[12] (Sprite_writeAddr[12]), .\Sprite_writeAddr[13] (Sprite_writeAddr[13]), 
            .\Sprite_readAddr[10] (Sprite_readAddr[10]), .Sprite_readData({Sprite_readData})) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    LUT_RAM RedLut (.\BUS_data[8] (BUS_data[8]), .\BUS_data[7] (BUS_data[7]), 
            .\BUS_data[6] (BUS_data[6]), .\BUS_data[5] (BUS_data[5]), .\BUS_data[4] (BUS_data[4]), 
            .\BUS_data[3] (BUS_data[3]), .\BUS_data[2] (BUS_data[2]), .\BUS_data[1] (BUS_data[1]), 
            .\BUS_data[0] (BUS_data[0]), .GND_net(GND_net), .\BUS_addr[10] (\BUS_addr[10] ), 
            .n17325(n17325), .n17337(n17337), .n17334(n17334), .n17321(n17321), 
            .n17331(n17331), .n17332(n17332), .n17333(n17333), .n17339(n17339), 
            .Sprite_readData({Sprite_readData}), .SpriteLut_writeClk(SpriteLut_writeClk), 
            .SpriteLut_readClk(SpriteLut_readClk), .VCC_net(VCC_net), .RED_WE(RED_WE), 
            .RED_WRITE({RED_WRITE}), .RED_READ({RED_READ})) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(651[11:18])
    LUT_RAM_U0 GreenLut (.\BUS_data[8] (BUS_data[8]), .\BUS_data[7] (BUS_data[7]), 
            .\BUS_data[6] (BUS_data[6]), .\BUS_data[5] (BUS_data[5]), .\BUS_data[4] (BUS_data[4]), 
            .\BUS_data[3] (BUS_data[3]), .\BUS_data[2] (BUS_data[2]), .\BUS_data[1] (BUS_data[1]), 
            .\BUS_data[0] (BUS_data[0]), .GND_net(GND_net), .\BUS_addr[10] (\BUS_addr[10] ), 
            .n17325(n17325), .n17337(n17337), .n17334(n17334), .n17321(n17321), 
            .n17331(n17331), .n17332(n17332), .n17333(n17333), .n17339(n17339), 
            .Sprite_readData({Sprite_readData}), .SpriteLut_writeClk(SpriteLut_writeClk), 
            .SpriteLut_readClk(SpriteLut_readClk), .VCC_net(VCC_net), .GREEN_WE(GREEN_WE), 
            .GREEN_WRITE({GREEN_WRITE}), .GREEN_READ({GREEN_READ})) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(669[12:19])
    GammaRam GRam (.\BUS_data[9] (BUS_data[9]), .GND_net(GND_net), .GR_WR_ADDR({GR_WR_ADDR}), 
            .currValue({currValue}), .GR_WR_CLK(GR_WR_CLK), .LOGIC_CLOCK_N_57(LOGIC_CLOCK_N_57), 
            .VCC_net(VCC_net), .n17387(n17387), .GR_WR_DOUT({GR_WR_DOUT}), 
            .GR_RE_DOUT({GR_RE_DOUT}), .\BUS_data[8] (BUS_data[8]), .\BUS_data[7] (BUS_data[7]), 
            .\BUS_data[6] (BUS_data[6]), .\BUS_data[5] (BUS_data[5]), .\BUS_data[4] (BUS_data[4]), 
            .\BUS_data[3] (BUS_data[3]), .\BUS_data[2] (BUS_data[2]), .\BUS_data[1] (BUS_data[1]), 
            .\BUS_data[0] (BUS_data[0])) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(616[8:16])
    LUT_RAM_U1 BlueLut (.\BUS_data[8] (BUS_data[8]), .\BUS_data[7] (BUS_data[7]), 
            .\BUS_data[6] (BUS_data[6]), .\BUS_data[5] (BUS_data[5]), .\BUS_data[4] (BUS_data[4]), 
            .\BUS_data[3] (BUS_data[3]), .\BUS_data[2] (BUS_data[2]), .\BUS_data[1] (BUS_data[1]), 
            .\BUS_data[0] (BUS_data[0]), .GND_net(GND_net), .\BUS_addr[10] (\BUS_addr[10] ), 
            .n17325(n17325), .n17337(n17337), .n17334(n17334), .n17321(n17321), 
            .n17331(n17331), .n17332(n17332), .n17333(n17333), .n17339(n17339), 
            .Sprite_readData({Sprite_readData}), .SpriteLut_writeClk(SpriteLut_writeClk), 
            .SpriteLut_readClk(SpriteLut_readClk), .VCC_net(VCC_net), .BLUE_WE(BLUE_WE), 
            .BLUE_WRITE({BLUE_WRITE}), .BLUE_READ({BLUE_READ})) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(687[11:18])
    LUT_RAM_U2 AlphaLut (.\BUS_data[8] (BUS_data[8]), .\BUS_data[7] (BUS_data[7]), 
            .\BUS_data[6] (BUS_data[6]), .\BUS_data[5] (BUS_data[5]), .\BUS_data[4] (BUS_data[4]), 
            .\BUS_data[3] (BUS_data[3]), .\BUS_data[2] (BUS_data[2]), .\BUS_data[1] (BUS_data[1]), 
            .\BUS_data[0] (BUS_data[0]), .GND_net(GND_net), .\BUS_addr[10] (\BUS_addr[10] ), 
            .n17325(n17325), .n17337(n17337), .n17334(n17334), .n17321(n17321), 
            .n17331(n17331), .n17332(n17332), .n17333(n17333), .n17339(n17339), 
            .Sprite_readData({Sprite_readData}), .SpriteLut_writeClk(SpriteLut_writeClk), 
            .SpriteLut_readClk(SpriteLut_readClk), .VCC_net(VCC_net), .ALPHA_WE(ALPHA_WE), 
            .ALPHA_WRITE({ALPHA_WRITE}), .ALPHA_READ({ALPHA_READ})) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(705[12:19])
    
endmodule
//
// Verilog Description of module SpriteRam
//

module SpriteRam (\Sprite_writeAddr[9] , \Sprite_writeAddr[8] , \Sprite_writeAddr[7] , 
            \Sprite_writeAddr[6] , \Sprite_writeAddr[5] , \Sprite_writeAddr[4] , 
            \Sprite_writeAddr[3] , \Sprite_writeAddr[2] , \Sprite_writeAddr[1] , 
            \Sprite_writeAddr[0] , \Sprite_readAddr[9] , \Sprite_readAddr[8] , 
            \Sprite_readAddr[7] , \Sprite_readAddr[6] , \Sprite_readAddr[5] , 
            \Sprite_readAddr[4] , \Sprite_readAddr[3] , \Sprite_readAddr[2] , 
            \Sprite_readAddr[1] , \Sprite_readAddr[0] , Sprite_writeData, 
            VCC_net, Sprite_readClk, GND_net, Sprite_writeClk, \Sprite_readAddr[11] , 
            \Sprite_readAddr[12] , \Sprite_readAddr[13] , \Sprite_writeAddr[11] , 
            \Sprite_writeAddr[10] , \Sprite_writeAddr[12] , \Sprite_writeAddr[13] , 
            \Sprite_readAddr[10] , Sprite_readData) /* synthesis NGD_DRC_MASK=1 */ ;
    input \Sprite_writeAddr[9] ;
    input \Sprite_writeAddr[8] ;
    input \Sprite_writeAddr[7] ;
    input \Sprite_writeAddr[6] ;
    input \Sprite_writeAddr[5] ;
    input \Sprite_writeAddr[4] ;
    input \Sprite_writeAddr[3] ;
    input \Sprite_writeAddr[2] ;
    input \Sprite_writeAddr[1] ;
    input \Sprite_writeAddr[0] ;
    input \Sprite_readAddr[9] ;
    input \Sprite_readAddr[8] ;
    input \Sprite_readAddr[7] ;
    input \Sprite_readAddr[6] ;
    input \Sprite_readAddr[5] ;
    input \Sprite_readAddr[4] ;
    input \Sprite_readAddr[3] ;
    input \Sprite_readAddr[2] ;
    input \Sprite_readAddr[1] ;
    input \Sprite_readAddr[0] ;
    input [8:0]Sprite_writeData;
    input VCC_net;
    input Sprite_readClk;
    input GND_net;
    input Sprite_writeClk;
    input \Sprite_readAddr[11] ;
    input \Sprite_readAddr[12] ;
    input \Sprite_readAddr[13] ;
    input \Sprite_writeAddr[11] ;
    input \Sprite_writeAddr[10] ;
    input \Sprite_writeAddr[12] ;
    input \Sprite_writeAddr[13] ;
    input \Sprite_readAddr[10] ;
    output [8:0]Sprite_readData;
    
    wire Sprite_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[9:23])
    wire Sprite_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(179[9:24])
    
    wire n15860, n15861, raddr11_ff, n15868, n15862, n15863, n15869, 
        mdout1_4_0, mdout1_5_0, raddr10_ff, n15864, n15865, n15870, 
        dec31_r115, dec30_p015, mdout1_15_0, mdout1_15_1, mdout1_15_2, 
        mdout1_15_3, mdout1_15_4, mdout1_15_5, mdout1_15_6, mdout1_15_7, 
        mdout1_15_8, n15866, n15867, n15871, raddr12_ff, raddr13_ff, 
        waddr11_inv, waddr10_inv, waddr12_inv, waddr13_inv, dec0_p00, 
        raddr10_inv, raddr11_inv, raddr12_inv, raddr13_inv, dec1_r10, 
        dec2_p01, dec3_r11, dec4_p02, dec5_r12, dec6_p03, dec7_r13, 
        dec8_p04, dec9_r14, dec10_p05, dec11_r15, dec12_p06, dec13_r16, 
        dec14_p07, dec15_r17, dec16_p08, dec17_r18, dec18_p09, dec19_r19, 
        dec20_p010, dec21_r110, dec22_p011, dec23_r111, dec24_p012, 
        dec25_r112, dec26_p013, dec27_r113, dec28_p014, dec29_r114, 
        mdout1_0_0, mdout1_0_1, mdout1_0_2, mdout1_0_3, mdout1_0_4, 
        mdout1_0_5, mdout1_0_6, mdout1_0_7, mdout1_0_8, mdout1_1_0, 
        mdout1_1_1, mdout1_1_2, mdout1_1_3, mdout1_1_4, mdout1_1_5, 
        mdout1_1_6, mdout1_1_7, mdout1_1_8, mdout1_2_0, mdout1_2_1, 
        mdout1_2_2, mdout1_2_3, mdout1_2_4, mdout1_2_5, mdout1_2_6, 
        mdout1_2_7, mdout1_2_8, mdout1_3_0, mdout1_3_1, mdout1_3_2, 
        mdout1_3_3, mdout1_3_4, mdout1_3_5, mdout1_3_6, mdout1_3_7, 
        mdout1_3_8, mdout1_4_1, mdout1_4_2, mdout1_4_3, mdout1_4_4, 
        mdout1_4_5, mdout1_4_6, mdout1_4_7, mdout1_4_8, mdout1_5_1, 
        mdout1_5_2, mdout1_5_3, mdout1_5_4, mdout1_5_5, mdout1_5_6, 
        mdout1_5_7, mdout1_5_8, mdout1_6_0, mdout1_6_1, mdout1_6_2, 
        mdout1_6_3, mdout1_6_4, mdout1_6_5, mdout1_6_6, mdout1_6_7, 
        mdout1_6_8, mdout1_7_0, mdout1_7_1, mdout1_7_2, mdout1_7_3, 
        mdout1_7_4, mdout1_7_5, mdout1_7_6, mdout1_7_7, mdout1_7_8, 
        mdout1_8_0, mdout1_8_1, mdout1_8_2, mdout1_8_3, mdout1_8_4, 
        mdout1_8_5, mdout1_8_6, mdout1_8_7, mdout1_8_8, mdout1_9_0, 
        mdout1_9_1, mdout1_9_2, mdout1_9_3, mdout1_9_4, mdout1_9_5, 
        mdout1_9_6, mdout1_9_7, mdout1_9_8, mdout1_10_0, mdout1_10_1, 
        mdout1_10_2, mdout1_10_3, mdout1_10_4, mdout1_10_5, mdout1_10_6, 
        mdout1_10_7, mdout1_10_8, mdout1_11_0, mdout1_11_1, mdout1_11_2, 
        mdout1_11_3, mdout1_11_4, mdout1_11_5, mdout1_11_6, mdout1_11_7, 
        mdout1_11_8, mdout1_12_0, mdout1_12_1, mdout1_12_2, mdout1_12_3, 
        mdout1_12_4, mdout1_12_5, mdout1_12_6, mdout1_12_7, mdout1_12_8, 
        mdout1_13_0, mdout1_13_1, mdout1_13_2, mdout1_13_3, mdout1_13_4, 
        mdout1_13_5, mdout1_13_6, mdout1_13_7, mdout1_13_8, mdout1_14_0, 
        mdout1_14_1, mdout1_14_2, mdout1_14_3, mdout1_14_4, mdout1_14_5, 
        mdout1_14_6, mdout1_14_7, mdout1_14_8, n15890, n15891, n15898, 
        n15880, n15879, n15897, n15896, n15987, n15878, n15986, 
        n15985, n15984, n15983, n15875, n15876, n15883, n15982, 
        n15981, n15980, n15972, n15971, n15970, n15969, n15968, 
        n15967, n15966, n15965, n15957, n15956, n15955, n15954, 
        n15953, n15952, n15951, n15950, n15942, n15941, n15940, 
        n15939, n15938, n15937, n15936, n15935, n15927, n15926, 
        n15925, n15924, n15923, n15922, n15921, n15920, n15912, 
        n15911, n15910, n15892, n15893, n15899, n15909, n15895, 
        n15908, n15907, n15906, n15905, n15894, n15877, n15884, 
        n15902, n15903, n15917, n15918, n15932, n15933, n15947, 
        n15948, n15962, n15963, n15977, n15978, n15992, n15993, 
        n15872, n15873, n15887, n15888, n15900, n15901, n15913, 
        n15914, n15915, n15916, n15928, n15929, n15930, n15931, 
        n15943, n15944, n15945, n15946, n15958, n15959, n15960, 
        n15961, n15973, n15974, n15975, n15976, n15988, n15989, 
        n15990, n15991, n15885, n15886, n15882, n15881;
    
    PFUMX i12206 (.BLUT(n15860), .ALUT(n15861), .C0(raddr11_ff), .Z(n15868));
    PFUMX i12207 (.BLUT(n15862), .ALUT(n15863), .C0(raddr11_ff), .Z(n15869));
    LUT4 i12200_3_lut (.A(mdout1_4_0), .B(mdout1_5_0), .C(raddr10_ff), 
         .Z(n15862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12200_3_lut.init = 16'hcaca;
    PFUMX i12208 (.BLUT(n15864), .ALUT(n15865), .C0(raddr11_ff), .Z(n15870));
    DP8KC SpriteRam_15_0_0 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec30_p015), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec31_r115), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_15_0), .DOB1(mdout1_15_1), 
          .DOB2(mdout1_15_2), .DOB3(mdout1_15_3), .DOB4(mdout1_15_4), 
          .DOB5(mdout1_15_5), .DOB6(mdout1_15_6), .DOB7(mdout1_15_7), 
          .DOB8(mdout1_15_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_15_0_0.DATA_WIDTH_A = 9;
    defparam SpriteRam_15_0_0.DATA_WIDTH_B = 9;
    defparam SpriteRam_15_0_0.REGMODE_A = "NOREG";
    defparam SpriteRam_15_0_0.REGMODE_B = "NOREG";
    defparam SpriteRam_15_0_0.CSDECODE_A = "0b001";
    defparam SpriteRam_15_0_0.CSDECODE_B = "0b001";
    defparam SpriteRam_15_0_0.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_15_0_0.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_15_0_0.GSR = "ENABLED";
    defparam SpriteRam_15_0_0.RESETMODE = "ASYNC";
    defparam SpriteRam_15_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_15_0_0.INIT_DATA = "STATIC";
    defparam SpriteRam_15_0_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_15_0_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PFUMX i12209 (.BLUT(n15866), .ALUT(n15867), .C0(raddr11_ff), .Z(n15871));
    FD1P3DX FF_2 (.D(\Sprite_readAddr[11] ), .SP(VCC_net), .CK(Sprite_readClk), 
            .CD(GND_net), .Q(raddr11_ff)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/spriteram.vhd(1554[11:18])
    defparam FF_2.GSR = "DISABLED";
    FD1P3DX FF_1 (.D(\Sprite_readAddr[12] ), .SP(VCC_net), .CK(Sprite_readClk), 
            .CD(GND_net), .Q(raddr12_ff)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/spriteram.vhd(1558[11:18])
    defparam FF_1.GSR = "DISABLED";
    FD1P3DX FF_0 (.D(\Sprite_readAddr[13] ), .SP(VCC_net), .CK(Sprite_readClk), 
            .CD(GND_net), .Q(raddr13_ff)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/spriteram.vhd(1565[11:18])
    defparam FF_0.GSR = "DISABLED";
    INV INV_6 (.A(\Sprite_writeAddr[11] ), .Z(waddr11_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    INV INV_7 (.A(\Sprite_writeAddr[10] ), .Z(waddr10_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    INV INV_5 (.A(\Sprite_writeAddr[12] ), .Z(waddr12_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    INV INV_4 (.A(\Sprite_writeAddr[13] ), .Z(waddr13_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    ROM16X1A LUT4_31 (.AD0(waddr13_inv), .AD1(waddr12_inv), .AD2(waddr11_inv), 
            .AD3(waddr10_inv), .DO0(dec0_p00)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_31.initval = 16'b1000000000000000;
    INV INV_3 (.A(\Sprite_readAddr[10] ), .Z(raddr10_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    INV INV_2 (.A(\Sprite_readAddr[11] ), .Z(raddr11_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    INV INV_1 (.A(\Sprite_readAddr[12] ), .Z(raddr12_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    INV INV_0 (.A(\Sprite_readAddr[13] ), .Z(raddr13_inv)) /* synthesis LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    ROM16X1A LUT4_30 (.AD0(raddr13_inv), .AD1(raddr12_inv), .AD2(raddr11_inv), 
            .AD3(raddr10_inv), .DO0(dec1_r10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_30.initval = 16'b1000000000000000;
    ROM16X1A LUT4_29 (.AD0(waddr13_inv), .AD1(waddr12_inv), .AD2(waddr11_inv), 
            .AD3(\Sprite_writeAddr[10] ), .DO0(dec2_p01)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_29.initval = 16'b1000000000000000;
    ROM16X1A LUT4_28 (.AD0(raddr13_inv), .AD1(raddr12_inv), .AD2(raddr11_inv), 
            .AD3(\Sprite_readAddr[10] ), .DO0(dec3_r11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_28.initval = 16'b1000000000000000;
    ROM16X1A LUT4_27 (.AD0(waddr13_inv), .AD1(waddr12_inv), .AD2(\Sprite_writeAddr[11] ), 
            .AD3(waddr10_inv), .DO0(dec4_p02)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_27.initval = 16'b1000000000000000;
    ROM16X1A LUT4_26 (.AD0(raddr13_inv), .AD1(raddr12_inv), .AD2(\Sprite_readAddr[11] ), 
            .AD3(raddr10_inv), .DO0(dec5_r12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_26.initval = 16'b1000000000000000;
    ROM16X1A LUT4_25 (.AD0(waddr13_inv), .AD1(waddr12_inv), .AD2(\Sprite_writeAddr[11] ), 
            .AD3(\Sprite_writeAddr[10] ), .DO0(dec6_p03)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_25.initval = 16'b1000000000000000;
    ROM16X1A LUT4_24 (.AD0(raddr13_inv), .AD1(raddr12_inv), .AD2(\Sprite_readAddr[11] ), 
            .AD3(\Sprite_readAddr[10] ), .DO0(dec7_r13)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_24.initval = 16'b1000000000000000;
    ROM16X1A LUT4_23 (.AD0(waddr13_inv), .AD1(\Sprite_writeAddr[12] ), .AD2(waddr11_inv), 
            .AD3(waddr10_inv), .DO0(dec8_p04)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_23.initval = 16'b1000000000000000;
    ROM16X1A LUT4_22 (.AD0(raddr13_inv), .AD1(\Sprite_readAddr[12] ), .AD2(raddr11_inv), 
            .AD3(raddr10_inv), .DO0(dec9_r14)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_22.initval = 16'b1000000000000000;
    ROM16X1A LUT4_21 (.AD0(waddr13_inv), .AD1(\Sprite_writeAddr[12] ), .AD2(waddr11_inv), 
            .AD3(\Sprite_writeAddr[10] ), .DO0(dec10_p05)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_21.initval = 16'b1000000000000000;
    ROM16X1A LUT4_20 (.AD0(raddr13_inv), .AD1(\Sprite_readAddr[12] ), .AD2(raddr11_inv), 
            .AD3(\Sprite_readAddr[10] ), .DO0(dec11_r15)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_20.initval = 16'b1000000000000000;
    ROM16X1A LUT4_19 (.AD0(waddr13_inv), .AD1(\Sprite_writeAddr[12] ), .AD2(\Sprite_writeAddr[11] ), 
            .AD3(waddr10_inv), .DO0(dec12_p06)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_19.initval = 16'b1000000000000000;
    ROM16X1A LUT4_18 (.AD0(raddr13_inv), .AD1(\Sprite_readAddr[12] ), .AD2(\Sprite_readAddr[11] ), 
            .AD3(raddr10_inv), .DO0(dec13_r16)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_18.initval = 16'b1000000000000000;
    ROM16X1A LUT4_17 (.AD0(waddr13_inv), .AD1(\Sprite_writeAddr[12] ), .AD2(\Sprite_writeAddr[11] ), 
            .AD3(\Sprite_writeAddr[10] ), .DO0(dec14_p07)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_17.initval = 16'b1000000000000000;
    ROM16X1A LUT4_16 (.AD0(raddr13_inv), .AD1(\Sprite_readAddr[12] ), .AD2(\Sprite_readAddr[11] ), 
            .AD3(\Sprite_readAddr[10] ), .DO0(dec15_r17)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_16.initval = 16'b1000000000000000;
    ROM16X1A LUT4_15 (.AD0(\Sprite_writeAddr[13] ), .AD1(waddr12_inv), .AD2(waddr11_inv), 
            .AD3(waddr10_inv), .DO0(dec16_p08)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_15.initval = 16'b1000000000000000;
    ROM16X1A LUT4_14 (.AD0(\Sprite_readAddr[13] ), .AD1(raddr12_inv), .AD2(raddr11_inv), 
            .AD3(raddr10_inv), .DO0(dec17_r18)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_14.initval = 16'b1000000000000000;
    ROM16X1A LUT4_13 (.AD0(\Sprite_writeAddr[13] ), .AD1(waddr12_inv), .AD2(waddr11_inv), 
            .AD3(\Sprite_writeAddr[10] ), .DO0(dec18_p09)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_13.initval = 16'b1000000000000000;
    ROM16X1A LUT4_12 (.AD0(\Sprite_readAddr[13] ), .AD1(raddr12_inv), .AD2(raddr11_inv), 
            .AD3(\Sprite_readAddr[10] ), .DO0(dec19_r19)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_12.initval = 16'b1000000000000000;
    ROM16X1A LUT4_11 (.AD0(\Sprite_writeAddr[13] ), .AD1(waddr12_inv), .AD2(\Sprite_writeAddr[11] ), 
            .AD3(waddr10_inv), .DO0(dec20_p010)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_11.initval = 16'b1000000000000000;
    ROM16X1A LUT4_10 (.AD0(\Sprite_readAddr[13] ), .AD1(raddr12_inv), .AD2(\Sprite_readAddr[11] ), 
            .AD3(raddr10_inv), .DO0(dec21_r110)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_10.initval = 16'b1000000000000000;
    ROM16X1A LUT4_9 (.AD0(\Sprite_writeAddr[13] ), .AD1(waddr12_inv), .AD2(\Sprite_writeAddr[11] ), 
            .AD3(\Sprite_writeAddr[10] ), .DO0(dec22_p011)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_9.initval = 16'b1000000000000000;
    ROM16X1A LUT4_8 (.AD0(\Sprite_readAddr[13] ), .AD1(raddr12_inv), .AD2(\Sprite_readAddr[11] ), 
            .AD3(\Sprite_readAddr[10] ), .DO0(dec23_r111)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_8.initval = 16'b1000000000000000;
    ROM16X1A LUT4_7 (.AD0(\Sprite_writeAddr[13] ), .AD1(\Sprite_writeAddr[12] ), 
            .AD2(waddr11_inv), .AD3(waddr10_inv), .DO0(dec24_p012)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_7.initval = 16'b1000000000000000;
    ROM16X1A LUT4_6 (.AD0(\Sprite_readAddr[13] ), .AD1(\Sprite_readAddr[12] ), 
            .AD2(raddr11_inv), .AD3(raddr10_inv), .DO0(dec25_r112)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_6.initval = 16'b1000000000000000;
    ROM16X1A LUT4_5 (.AD0(\Sprite_writeAddr[13] ), .AD1(\Sprite_writeAddr[12] ), 
            .AD2(waddr11_inv), .AD3(\Sprite_writeAddr[10] ), .DO0(dec26_p013)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_5.initval = 16'b1000000000000000;
    ROM16X1A LUT4_4 (.AD0(\Sprite_readAddr[13] ), .AD1(\Sprite_readAddr[12] ), 
            .AD2(raddr11_inv), .AD3(\Sprite_readAddr[10] ), .DO0(dec27_r113)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_4.initval = 16'b1000000000000000;
    ROM16X1A LUT4_3 (.AD0(\Sprite_writeAddr[13] ), .AD1(\Sprite_writeAddr[12] ), 
            .AD2(\Sprite_writeAddr[11] ), .AD3(waddr10_inv), .DO0(dec28_p014)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_3.initval = 16'b1000000000000000;
    ROM16X1A LUT4_2 (.AD0(\Sprite_readAddr[13] ), .AD1(\Sprite_readAddr[12] ), 
            .AD2(\Sprite_readAddr[11] ), .AD3(raddr10_inv), .DO0(dec29_r114)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_2.initval = 16'b1000000000000000;
    ROM16X1A LUT4_1 (.AD0(\Sprite_writeAddr[13] ), .AD1(\Sprite_writeAddr[12] ), 
            .AD2(\Sprite_writeAddr[11] ), .AD3(\Sprite_writeAddr[10] ), 
            .DO0(dec30_p015)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_1.initval = 16'b1000000000000000;
    ROM16X1A LUT4_0 (.AD0(\Sprite_readAddr[13] ), .AD1(\Sprite_readAddr[12] ), 
            .AD2(\Sprite_readAddr[11] ), .AD3(\Sprite_readAddr[10] ), .DO0(dec31_r115)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam LUT4_0.initval = 16'b1000000000000000;
    DP8KC SpriteRam_0_0_15 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec0_p00), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec1_r10), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_0_0), .DOB1(mdout1_0_1), 
          .DOB2(mdout1_0_2), .DOB3(mdout1_0_3), .DOB4(mdout1_0_4), .DOB5(mdout1_0_5), 
          .DOB6(mdout1_0_6), .DOB7(mdout1_0_7), .DOB8(mdout1_0_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_0_0_15.DATA_WIDTH_A = 9;
    defparam SpriteRam_0_0_15.DATA_WIDTH_B = 9;
    defparam SpriteRam_0_0_15.REGMODE_A = "NOREG";
    defparam SpriteRam_0_0_15.REGMODE_B = "NOREG";
    defparam SpriteRam_0_0_15.CSDECODE_A = "0b001";
    defparam SpriteRam_0_0_15.CSDECODE_B = "0b001";
    defparam SpriteRam_0_0_15.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_0_0_15.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_0_0_15.GSR = "ENABLED";
    defparam SpriteRam_0_0_15.RESETMODE = "ASYNC";
    defparam SpriteRam_0_0_15.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_0_0_15.INIT_DATA = "STATIC";
    defparam SpriteRam_0_0_15.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_0_0_15.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_1_0_14 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec2_p01), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec3_r11), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_1_0), .DOB1(mdout1_1_1), 
          .DOB2(mdout1_1_2), .DOB3(mdout1_1_3), .DOB4(mdout1_1_4), .DOB5(mdout1_1_5), 
          .DOB6(mdout1_1_6), .DOB7(mdout1_1_7), .DOB8(mdout1_1_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_1_0_14.DATA_WIDTH_A = 9;
    defparam SpriteRam_1_0_14.DATA_WIDTH_B = 9;
    defparam SpriteRam_1_0_14.REGMODE_A = "NOREG";
    defparam SpriteRam_1_0_14.REGMODE_B = "NOREG";
    defparam SpriteRam_1_0_14.CSDECODE_A = "0b001";
    defparam SpriteRam_1_0_14.CSDECODE_B = "0b001";
    defparam SpriteRam_1_0_14.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_1_0_14.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_1_0_14.GSR = "ENABLED";
    defparam SpriteRam_1_0_14.RESETMODE = "ASYNC";
    defparam SpriteRam_1_0_14.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_1_0_14.INIT_DATA = "STATIC";
    defparam SpriteRam_1_0_14.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_1_0_14.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_2_0_13 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec4_p02), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec5_r12), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_2_0), .DOB1(mdout1_2_1), 
          .DOB2(mdout1_2_2), .DOB3(mdout1_2_3), .DOB4(mdout1_2_4), .DOB5(mdout1_2_5), 
          .DOB6(mdout1_2_6), .DOB7(mdout1_2_7), .DOB8(mdout1_2_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_2_0_13.DATA_WIDTH_A = 9;
    defparam SpriteRam_2_0_13.DATA_WIDTH_B = 9;
    defparam SpriteRam_2_0_13.REGMODE_A = "NOREG";
    defparam SpriteRam_2_0_13.REGMODE_B = "NOREG";
    defparam SpriteRam_2_0_13.CSDECODE_A = "0b001";
    defparam SpriteRam_2_0_13.CSDECODE_B = "0b001";
    defparam SpriteRam_2_0_13.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_2_0_13.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_2_0_13.GSR = "ENABLED";
    defparam SpriteRam_2_0_13.RESETMODE = "ASYNC";
    defparam SpriteRam_2_0_13.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_2_0_13.INIT_DATA = "STATIC";
    defparam SpriteRam_2_0_13.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_2_0_13.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_3_0_12 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec6_p03), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec7_r13), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_3_0), .DOB1(mdout1_3_1), 
          .DOB2(mdout1_3_2), .DOB3(mdout1_3_3), .DOB4(mdout1_3_4), .DOB5(mdout1_3_5), 
          .DOB6(mdout1_3_6), .DOB7(mdout1_3_7), .DOB8(mdout1_3_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_3_0_12.DATA_WIDTH_A = 9;
    defparam SpriteRam_3_0_12.DATA_WIDTH_B = 9;
    defparam SpriteRam_3_0_12.REGMODE_A = "NOREG";
    defparam SpriteRam_3_0_12.REGMODE_B = "NOREG";
    defparam SpriteRam_3_0_12.CSDECODE_A = "0b001";
    defparam SpriteRam_3_0_12.CSDECODE_B = "0b001";
    defparam SpriteRam_3_0_12.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_3_0_12.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_3_0_12.GSR = "ENABLED";
    defparam SpriteRam_3_0_12.RESETMODE = "ASYNC";
    defparam SpriteRam_3_0_12.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_3_0_12.INIT_DATA = "STATIC";
    defparam SpriteRam_3_0_12.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_3_0_12.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_4_0_11 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec8_p04), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec9_r14), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_4_0), .DOB1(mdout1_4_1), 
          .DOB2(mdout1_4_2), .DOB3(mdout1_4_3), .DOB4(mdout1_4_4), .DOB5(mdout1_4_5), 
          .DOB6(mdout1_4_6), .DOB7(mdout1_4_7), .DOB8(mdout1_4_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_4_0_11.DATA_WIDTH_A = 9;
    defparam SpriteRam_4_0_11.DATA_WIDTH_B = 9;
    defparam SpriteRam_4_0_11.REGMODE_A = "NOREG";
    defparam SpriteRam_4_0_11.REGMODE_B = "NOREG";
    defparam SpriteRam_4_0_11.CSDECODE_A = "0b001";
    defparam SpriteRam_4_0_11.CSDECODE_B = "0b001";
    defparam SpriteRam_4_0_11.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_4_0_11.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_4_0_11.GSR = "ENABLED";
    defparam SpriteRam_4_0_11.RESETMODE = "ASYNC";
    defparam SpriteRam_4_0_11.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_4_0_11.INIT_DATA = "STATIC";
    defparam SpriteRam_4_0_11.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_4_0_11.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_5_0_10 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec10_p05), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec11_r15), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_5_0), .DOB1(mdout1_5_1), 
          .DOB2(mdout1_5_2), .DOB3(mdout1_5_3), .DOB4(mdout1_5_4), .DOB5(mdout1_5_5), 
          .DOB6(mdout1_5_6), .DOB7(mdout1_5_7), .DOB8(mdout1_5_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_5_0_10.DATA_WIDTH_A = 9;
    defparam SpriteRam_5_0_10.DATA_WIDTH_B = 9;
    defparam SpriteRam_5_0_10.REGMODE_A = "NOREG";
    defparam SpriteRam_5_0_10.REGMODE_B = "NOREG";
    defparam SpriteRam_5_0_10.CSDECODE_A = "0b001";
    defparam SpriteRam_5_0_10.CSDECODE_B = "0b001";
    defparam SpriteRam_5_0_10.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_5_0_10.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_5_0_10.GSR = "ENABLED";
    defparam SpriteRam_5_0_10.RESETMODE = "ASYNC";
    defparam SpriteRam_5_0_10.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_5_0_10.INIT_DATA = "STATIC";
    defparam SpriteRam_5_0_10.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_5_0_10.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_6_0_9 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec12_p06), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec13_r16), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_6_0), .DOB1(mdout1_6_1), 
          .DOB2(mdout1_6_2), .DOB3(mdout1_6_3), .DOB4(mdout1_6_4), .DOB5(mdout1_6_5), 
          .DOB6(mdout1_6_6), .DOB7(mdout1_6_7), .DOB8(mdout1_6_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_6_0_9.DATA_WIDTH_A = 9;
    defparam SpriteRam_6_0_9.DATA_WIDTH_B = 9;
    defparam SpriteRam_6_0_9.REGMODE_A = "NOREG";
    defparam SpriteRam_6_0_9.REGMODE_B = "NOREG";
    defparam SpriteRam_6_0_9.CSDECODE_A = "0b001";
    defparam SpriteRam_6_0_9.CSDECODE_B = "0b001";
    defparam SpriteRam_6_0_9.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_6_0_9.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_6_0_9.GSR = "ENABLED";
    defparam SpriteRam_6_0_9.RESETMODE = "ASYNC";
    defparam SpriteRam_6_0_9.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_6_0_9.INIT_DATA = "STATIC";
    defparam SpriteRam_6_0_9.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_6_0_9.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_7_0_8 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec14_p07), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec15_r17), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_7_0), .DOB1(mdout1_7_1), 
          .DOB2(mdout1_7_2), .DOB3(mdout1_7_3), .DOB4(mdout1_7_4), .DOB5(mdout1_7_5), 
          .DOB6(mdout1_7_6), .DOB7(mdout1_7_7), .DOB8(mdout1_7_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_7_0_8.DATA_WIDTH_A = 9;
    defparam SpriteRam_7_0_8.DATA_WIDTH_B = 9;
    defparam SpriteRam_7_0_8.REGMODE_A = "NOREG";
    defparam SpriteRam_7_0_8.REGMODE_B = "NOREG";
    defparam SpriteRam_7_0_8.CSDECODE_A = "0b001";
    defparam SpriteRam_7_0_8.CSDECODE_B = "0b001";
    defparam SpriteRam_7_0_8.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_7_0_8.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_7_0_8.GSR = "ENABLED";
    defparam SpriteRam_7_0_8.RESETMODE = "ASYNC";
    defparam SpriteRam_7_0_8.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_7_0_8.INIT_DATA = "STATIC";
    defparam SpriteRam_7_0_8.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_7_0_8.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_8_0_7 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec16_p08), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec17_r18), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_8_0), .DOB1(mdout1_8_1), 
          .DOB2(mdout1_8_2), .DOB3(mdout1_8_3), .DOB4(mdout1_8_4), .DOB5(mdout1_8_5), 
          .DOB6(mdout1_8_6), .DOB7(mdout1_8_7), .DOB8(mdout1_8_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_8_0_7.DATA_WIDTH_A = 9;
    defparam SpriteRam_8_0_7.DATA_WIDTH_B = 9;
    defparam SpriteRam_8_0_7.REGMODE_A = "NOREG";
    defparam SpriteRam_8_0_7.REGMODE_B = "NOREG";
    defparam SpriteRam_8_0_7.CSDECODE_A = "0b001";
    defparam SpriteRam_8_0_7.CSDECODE_B = "0b001";
    defparam SpriteRam_8_0_7.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_8_0_7.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_8_0_7.GSR = "ENABLED";
    defparam SpriteRam_8_0_7.RESETMODE = "ASYNC";
    defparam SpriteRam_8_0_7.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_8_0_7.INIT_DATA = "STATIC";
    defparam SpriteRam_8_0_7.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_8_0_7.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_9_0_6 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec18_p09), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec19_r19), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_9_0), .DOB1(mdout1_9_1), 
          .DOB2(mdout1_9_2), .DOB3(mdout1_9_3), .DOB4(mdout1_9_4), .DOB5(mdout1_9_5), 
          .DOB6(mdout1_9_6), .DOB7(mdout1_9_7), .DOB8(mdout1_9_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_9_0_6.DATA_WIDTH_A = 9;
    defparam SpriteRam_9_0_6.DATA_WIDTH_B = 9;
    defparam SpriteRam_9_0_6.REGMODE_A = "NOREG";
    defparam SpriteRam_9_0_6.REGMODE_B = "NOREG";
    defparam SpriteRam_9_0_6.CSDECODE_A = "0b001";
    defparam SpriteRam_9_0_6.CSDECODE_B = "0b001";
    defparam SpriteRam_9_0_6.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_9_0_6.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_9_0_6.GSR = "ENABLED";
    defparam SpriteRam_9_0_6.RESETMODE = "ASYNC";
    defparam SpriteRam_9_0_6.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_9_0_6.INIT_DATA = "STATIC";
    defparam SpriteRam_9_0_6.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_9_0_6.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_10_0_5 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec20_p010), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec21_r110), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_10_0), .DOB1(mdout1_10_1), 
          .DOB2(mdout1_10_2), .DOB3(mdout1_10_3), .DOB4(mdout1_10_4), 
          .DOB5(mdout1_10_5), .DOB6(mdout1_10_6), .DOB7(mdout1_10_7), 
          .DOB8(mdout1_10_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_10_0_5.DATA_WIDTH_A = 9;
    defparam SpriteRam_10_0_5.DATA_WIDTH_B = 9;
    defparam SpriteRam_10_0_5.REGMODE_A = "NOREG";
    defparam SpriteRam_10_0_5.REGMODE_B = "NOREG";
    defparam SpriteRam_10_0_5.CSDECODE_A = "0b001";
    defparam SpriteRam_10_0_5.CSDECODE_B = "0b001";
    defparam SpriteRam_10_0_5.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_10_0_5.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_10_0_5.GSR = "ENABLED";
    defparam SpriteRam_10_0_5.RESETMODE = "ASYNC";
    defparam SpriteRam_10_0_5.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_10_0_5.INIT_DATA = "STATIC";
    defparam SpriteRam_10_0_5.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_10_0_5.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_11_0_4 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec22_p011), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec23_r111), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_11_0), .DOB1(mdout1_11_1), 
          .DOB2(mdout1_11_2), .DOB3(mdout1_11_3), .DOB4(mdout1_11_4), 
          .DOB5(mdout1_11_5), .DOB6(mdout1_11_6), .DOB7(mdout1_11_7), 
          .DOB8(mdout1_11_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_11_0_4.DATA_WIDTH_A = 9;
    defparam SpriteRam_11_0_4.DATA_WIDTH_B = 9;
    defparam SpriteRam_11_0_4.REGMODE_A = "NOREG";
    defparam SpriteRam_11_0_4.REGMODE_B = "NOREG";
    defparam SpriteRam_11_0_4.CSDECODE_A = "0b001";
    defparam SpriteRam_11_0_4.CSDECODE_B = "0b001";
    defparam SpriteRam_11_0_4.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_11_0_4.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_11_0_4.GSR = "ENABLED";
    defparam SpriteRam_11_0_4.RESETMODE = "ASYNC";
    defparam SpriteRam_11_0_4.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_11_0_4.INIT_DATA = "STATIC";
    defparam SpriteRam_11_0_4.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_11_0_4.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_12_0_3 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec24_p012), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec25_r112), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_12_0), .DOB1(mdout1_12_1), 
          .DOB2(mdout1_12_2), .DOB3(mdout1_12_3), .DOB4(mdout1_12_4), 
          .DOB5(mdout1_12_5), .DOB6(mdout1_12_6), .DOB7(mdout1_12_7), 
          .DOB8(mdout1_12_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_12_0_3.DATA_WIDTH_A = 9;
    defparam SpriteRam_12_0_3.DATA_WIDTH_B = 9;
    defparam SpriteRam_12_0_3.REGMODE_A = "NOREG";
    defparam SpriteRam_12_0_3.REGMODE_B = "NOREG";
    defparam SpriteRam_12_0_3.CSDECODE_A = "0b001";
    defparam SpriteRam_12_0_3.CSDECODE_B = "0b001";
    defparam SpriteRam_12_0_3.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_12_0_3.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_12_0_3.GSR = "ENABLED";
    defparam SpriteRam_12_0_3.RESETMODE = "ASYNC";
    defparam SpriteRam_12_0_3.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_12_0_3.INIT_DATA = "STATIC";
    defparam SpriteRam_12_0_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_12_0_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_13_0_2 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec26_p013), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec27_r113), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_13_0), .DOB1(mdout1_13_1), 
          .DOB2(mdout1_13_2), .DOB3(mdout1_13_3), .DOB4(mdout1_13_4), 
          .DOB5(mdout1_13_5), .DOB6(mdout1_13_6), .DOB7(mdout1_13_7), 
          .DOB8(mdout1_13_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_13_0_2.DATA_WIDTH_A = 9;
    defparam SpriteRam_13_0_2.DATA_WIDTH_B = 9;
    defparam SpriteRam_13_0_2.REGMODE_A = "NOREG";
    defparam SpriteRam_13_0_2.REGMODE_B = "NOREG";
    defparam SpriteRam_13_0_2.CSDECODE_A = "0b001";
    defparam SpriteRam_13_0_2.CSDECODE_B = "0b001";
    defparam SpriteRam_13_0_2.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_13_0_2.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_13_0_2.GSR = "ENABLED";
    defparam SpriteRam_13_0_2.RESETMODE = "ASYNC";
    defparam SpriteRam_13_0_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_13_0_2.INIT_DATA = "STATIC";
    defparam SpriteRam_13_0_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_13_0_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC SpriteRam_14_0_1 (.DIA0(Sprite_writeData[0]), .DIA1(Sprite_writeData[1]), 
          .DIA2(Sprite_writeData[2]), .DIA3(Sprite_writeData[3]), .DIA4(Sprite_writeData[4]), 
          .DIA5(Sprite_writeData[5]), .DIA6(Sprite_writeData[6]), .DIA7(Sprite_writeData[7]), 
          .DIA8(Sprite_writeData[8]), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(\Sprite_writeAddr[0] ), .ADA4(\Sprite_writeAddr[1] ), 
          .ADA5(\Sprite_writeAddr[2] ), .ADA6(\Sprite_writeAddr[3] ), .ADA7(\Sprite_writeAddr[4] ), 
          .ADA8(\Sprite_writeAddr[5] ), .ADA9(\Sprite_writeAddr[6] ), .ADA10(\Sprite_writeAddr[7] ), 
          .ADA11(\Sprite_writeAddr[8] ), .ADA12(\Sprite_writeAddr[9] ), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(Sprite_writeClk), .WEA(VCC_net), 
          .CSA0(dec28_p014), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(\Sprite_readAddr[0] ), .ADB4(\Sprite_readAddr[1] ), .ADB5(\Sprite_readAddr[2] ), 
          .ADB6(\Sprite_readAddr[3] ), .ADB7(\Sprite_readAddr[4] ), .ADB8(\Sprite_readAddr[5] ), 
          .ADB9(\Sprite_readAddr[6] ), .ADB10(\Sprite_readAddr[7] ), .ADB11(\Sprite_readAddr[8] ), 
          .ADB12(\Sprite_readAddr[9] ), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(Sprite_readClk), .WEB(GND_net), .CSB0(dec29_r114), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOB0(mdout1_14_0), .DOB1(mdout1_14_1), 
          .DOB2(mdout1_14_2), .DOB3(mdout1_14_3), .DOB4(mdout1_14_4), 
          .DOB5(mdout1_14_5), .DOB6(mdout1_14_6), .DOB7(mdout1_14_7), 
          .DOB8(mdout1_14_8)) /* synthesis MEM_LPC_FILE="SpriteRam.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam SpriteRam_14_0_1.DATA_WIDTH_A = 9;
    defparam SpriteRam_14_0_1.DATA_WIDTH_B = 9;
    defparam SpriteRam_14_0_1.REGMODE_A = "NOREG";
    defparam SpriteRam_14_0_1.REGMODE_B = "NOREG";
    defparam SpriteRam_14_0_1.CSDECODE_A = "0b001";
    defparam SpriteRam_14_0_1.CSDECODE_B = "0b001";
    defparam SpriteRam_14_0_1.WRITEMODE_A = "NORMAL";
    defparam SpriteRam_14_0_1.WRITEMODE_B = "NORMAL";
    defparam SpriteRam_14_0_1.GSR = "ENABLED";
    defparam SpriteRam_14_0_1.RESETMODE = "ASYNC";
    defparam SpriteRam_14_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam SpriteRam_14_0_1.INIT_DATA = "STATIC";
    defparam SpriteRam_14_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam SpriteRam_14_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    FD1P3DX FF_3 (.D(\Sprite_readAddr[10] ), .SP(VCC_net), .CK(Sprite_readClk), 
            .CD(GND_net), .Q(raddr10_ff)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=17, LSE_LLINE=634, LSE_RLINE=634 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/spriteram.vhd(1550[11:18])
    defparam FF_3.GSR = "DISABLED";
    PFUMX i12236 (.BLUT(n15890), .ALUT(n15891), .C0(raddr11_ff), .Z(n15898));
    LUT4 i12218_3_lut (.A(mdout1_10_1), .B(mdout1_11_1), .C(raddr10_ff), 
         .Z(n15880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12218_3_lut.init = 16'hcaca;
    LUT4 i12217_3_lut (.A(mdout1_8_1), .B(mdout1_9_1), .C(raddr10_ff), 
         .Z(n15879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12217_3_lut.init = 16'hcaca;
    LUT4 i12235_3_lut (.A(mdout1_14_2), .B(mdout1_15_2), .C(raddr10_ff), 
         .Z(n15897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12235_3_lut.init = 16'hcaca;
    LUT4 i12234_3_lut (.A(mdout1_12_2), .B(mdout1_13_2), .C(raddr10_ff), 
         .Z(n15896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12234_3_lut.init = 16'hcaca;
    LUT4 i12325_3_lut (.A(mdout1_14_8), .B(mdout1_15_8), .C(raddr10_ff), 
         .Z(n15987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12325_3_lut.init = 16'hcaca;
    LUT4 i12216_3_lut (.A(mdout1_6_1), .B(mdout1_7_1), .C(raddr10_ff), 
         .Z(n15878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12216_3_lut.init = 16'hcaca;
    LUT4 i12324_3_lut (.A(mdout1_12_8), .B(mdout1_13_8), .C(raddr10_ff), 
         .Z(n15986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12324_3_lut.init = 16'hcaca;
    LUT4 i12323_3_lut (.A(mdout1_10_8), .B(mdout1_11_8), .C(raddr10_ff), 
         .Z(n15985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12323_3_lut.init = 16'hcaca;
    LUT4 i12322_3_lut (.A(mdout1_8_8), .B(mdout1_9_8), .C(raddr10_ff), 
         .Z(n15984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12322_3_lut.init = 16'hcaca;
    LUT4 i12321_3_lut (.A(mdout1_6_8), .B(mdout1_7_8), .C(raddr10_ff), 
         .Z(n15983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12321_3_lut.init = 16'hcaca;
    PFUMX i12221 (.BLUT(n15875), .ALUT(n15876), .C0(raddr11_ff), .Z(n15883));
    LUT4 i12320_3_lut (.A(mdout1_4_8), .B(mdout1_5_8), .C(raddr10_ff), 
         .Z(n15982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12320_3_lut.init = 16'hcaca;
    LUT4 i12319_3_lut (.A(mdout1_2_8), .B(mdout1_3_8), .C(raddr10_ff), 
         .Z(n15981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12319_3_lut.init = 16'hcaca;
    LUT4 i12318_3_lut (.A(mdout1_0_8), .B(mdout1_1_8), .C(raddr10_ff), 
         .Z(n15980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12318_3_lut.init = 16'hcaca;
    LUT4 i12310_3_lut (.A(mdout1_14_7), .B(mdout1_15_7), .C(raddr10_ff), 
         .Z(n15972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12310_3_lut.init = 16'hcaca;
    LUT4 i12309_3_lut (.A(mdout1_12_7), .B(mdout1_13_7), .C(raddr10_ff), 
         .Z(n15971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12309_3_lut.init = 16'hcaca;
    LUT4 i12308_3_lut (.A(mdout1_10_7), .B(mdout1_11_7), .C(raddr10_ff), 
         .Z(n15970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12308_3_lut.init = 16'hcaca;
    LUT4 i12307_3_lut (.A(mdout1_8_7), .B(mdout1_9_7), .C(raddr10_ff), 
         .Z(n15969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12307_3_lut.init = 16'hcaca;
    LUT4 i12306_3_lut (.A(mdout1_6_7), .B(mdout1_7_7), .C(raddr10_ff), 
         .Z(n15968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12306_3_lut.init = 16'hcaca;
    LUT4 i12305_3_lut (.A(mdout1_4_7), .B(mdout1_5_7), .C(raddr10_ff), 
         .Z(n15967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12305_3_lut.init = 16'hcaca;
    LUT4 i12304_3_lut (.A(mdout1_2_7), .B(mdout1_3_7), .C(raddr10_ff), 
         .Z(n15966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12304_3_lut.init = 16'hcaca;
    LUT4 i12303_3_lut (.A(mdout1_0_7), .B(mdout1_1_7), .C(raddr10_ff), 
         .Z(n15965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12303_3_lut.init = 16'hcaca;
    LUT4 i12295_3_lut (.A(mdout1_14_6), .B(mdout1_15_6), .C(raddr10_ff), 
         .Z(n15957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12295_3_lut.init = 16'hcaca;
    LUT4 i12294_3_lut (.A(mdout1_12_6), .B(mdout1_13_6), .C(raddr10_ff), 
         .Z(n15956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12294_3_lut.init = 16'hcaca;
    LUT4 i12293_3_lut (.A(mdout1_10_6), .B(mdout1_11_6), .C(raddr10_ff), 
         .Z(n15955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12293_3_lut.init = 16'hcaca;
    LUT4 i12292_3_lut (.A(mdout1_8_6), .B(mdout1_9_6), .C(raddr10_ff), 
         .Z(n15954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12292_3_lut.init = 16'hcaca;
    LUT4 i12291_3_lut (.A(mdout1_6_6), .B(mdout1_7_6), .C(raddr10_ff), 
         .Z(n15953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12291_3_lut.init = 16'hcaca;
    LUT4 i12290_3_lut (.A(mdout1_4_6), .B(mdout1_5_6), .C(raddr10_ff), 
         .Z(n15952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12290_3_lut.init = 16'hcaca;
    LUT4 i12289_3_lut (.A(mdout1_2_6), .B(mdout1_3_6), .C(raddr10_ff), 
         .Z(n15951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12289_3_lut.init = 16'hcaca;
    LUT4 i12288_3_lut (.A(mdout1_0_6), .B(mdout1_1_6), .C(raddr10_ff), 
         .Z(n15950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12288_3_lut.init = 16'hcaca;
    LUT4 i12280_3_lut (.A(mdout1_14_5), .B(mdout1_15_5), .C(raddr10_ff), 
         .Z(n15942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12280_3_lut.init = 16'hcaca;
    LUT4 i12279_3_lut (.A(mdout1_12_5), .B(mdout1_13_5), .C(raddr10_ff), 
         .Z(n15941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12279_3_lut.init = 16'hcaca;
    LUT4 i12278_3_lut (.A(mdout1_10_5), .B(mdout1_11_5), .C(raddr10_ff), 
         .Z(n15940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12278_3_lut.init = 16'hcaca;
    LUT4 i12277_3_lut (.A(mdout1_8_5), .B(mdout1_9_5), .C(raddr10_ff), 
         .Z(n15939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12277_3_lut.init = 16'hcaca;
    LUT4 i12276_3_lut (.A(mdout1_6_5), .B(mdout1_7_5), .C(raddr10_ff), 
         .Z(n15938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12276_3_lut.init = 16'hcaca;
    LUT4 i12275_3_lut (.A(mdout1_4_5), .B(mdout1_5_5), .C(raddr10_ff), 
         .Z(n15937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12275_3_lut.init = 16'hcaca;
    LUT4 i12274_3_lut (.A(mdout1_2_5), .B(mdout1_3_5), .C(raddr10_ff), 
         .Z(n15936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12274_3_lut.init = 16'hcaca;
    LUT4 i12273_3_lut (.A(mdout1_0_5), .B(mdout1_1_5), .C(raddr10_ff), 
         .Z(n15935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12273_3_lut.init = 16'hcaca;
    LUT4 i12265_3_lut (.A(mdout1_14_4), .B(mdout1_15_4), .C(raddr10_ff), 
         .Z(n15927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12265_3_lut.init = 16'hcaca;
    LUT4 i12264_3_lut (.A(mdout1_12_4), .B(mdout1_13_4), .C(raddr10_ff), 
         .Z(n15926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12264_3_lut.init = 16'hcaca;
    LUT4 i12263_3_lut (.A(mdout1_10_4), .B(mdout1_11_4), .C(raddr10_ff), 
         .Z(n15925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12263_3_lut.init = 16'hcaca;
    LUT4 i12262_3_lut (.A(mdout1_8_4), .B(mdout1_9_4), .C(raddr10_ff), 
         .Z(n15924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12262_3_lut.init = 16'hcaca;
    LUT4 i12261_3_lut (.A(mdout1_6_4), .B(mdout1_7_4), .C(raddr10_ff), 
         .Z(n15923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12261_3_lut.init = 16'hcaca;
    LUT4 i12260_3_lut (.A(mdout1_4_4), .B(mdout1_5_4), .C(raddr10_ff), 
         .Z(n15922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12260_3_lut.init = 16'hcaca;
    LUT4 i12259_3_lut (.A(mdout1_2_4), .B(mdout1_3_4), .C(raddr10_ff), 
         .Z(n15921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12259_3_lut.init = 16'hcaca;
    LUT4 i12258_3_lut (.A(mdout1_0_4), .B(mdout1_1_4), .C(raddr10_ff), 
         .Z(n15920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12258_3_lut.init = 16'hcaca;
    LUT4 i12250_3_lut (.A(mdout1_14_3), .B(mdout1_15_3), .C(raddr10_ff), 
         .Z(n15912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12250_3_lut.init = 16'hcaca;
    LUT4 i12249_3_lut (.A(mdout1_12_3), .B(mdout1_13_3), .C(raddr10_ff), 
         .Z(n15911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12249_3_lut.init = 16'hcaca;
    LUT4 i12248_3_lut (.A(mdout1_10_3), .B(mdout1_11_3), .C(raddr10_ff), 
         .Z(n15910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12248_3_lut.init = 16'hcaca;
    PFUMX i12237 (.BLUT(n15892), .ALUT(n15893), .C0(raddr11_ff), .Z(n15899));
    LUT4 i12247_3_lut (.A(mdout1_8_3), .B(mdout1_9_3), .C(raddr10_ff), 
         .Z(n15909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12247_3_lut.init = 16'hcaca;
    LUT4 i12233_3_lut (.A(mdout1_10_2), .B(mdout1_11_2), .C(raddr10_ff), 
         .Z(n15895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12233_3_lut.init = 16'hcaca;
    LUT4 i12246_3_lut (.A(mdout1_6_3), .B(mdout1_7_3), .C(raddr10_ff), 
         .Z(n15908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12246_3_lut.init = 16'hcaca;
    LUT4 i12245_3_lut (.A(mdout1_4_3), .B(mdout1_5_3), .C(raddr10_ff), 
         .Z(n15907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12245_3_lut.init = 16'hcaca;
    LUT4 i12244_3_lut (.A(mdout1_2_3), .B(mdout1_3_3), .C(raddr10_ff), 
         .Z(n15906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12244_3_lut.init = 16'hcaca;
    LUT4 i12243_3_lut (.A(mdout1_0_3), .B(mdout1_1_3), .C(raddr10_ff), 
         .Z(n15905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12243_3_lut.init = 16'hcaca;
    LUT4 i12232_3_lut (.A(mdout1_8_2), .B(mdout1_9_2), .C(raddr10_ff), 
         .Z(n15894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12232_3_lut.init = 16'hcaca;
    LUT4 i12231_3_lut (.A(mdout1_6_2), .B(mdout1_7_2), .C(raddr10_ff), 
         .Z(n15893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12231_3_lut.init = 16'hcaca;
    LUT4 i12230_3_lut (.A(mdout1_4_2), .B(mdout1_5_2), .C(raddr10_ff), 
         .Z(n15892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12230_3_lut.init = 16'hcaca;
    PFUMX i12222 (.BLUT(n15877), .ALUT(n15878), .C0(raddr11_ff), .Z(n15884));
    L6MUX21 i12242 (.D0(n15902), .D1(n15903), .SD(raddr13_ff), .Z(Sprite_readData[2]));
    L6MUX21 i12257 (.D0(n15917), .D1(n15918), .SD(raddr13_ff), .Z(Sprite_readData[3]));
    L6MUX21 i12272 (.D0(n15932), .D1(n15933), .SD(raddr13_ff), .Z(Sprite_readData[4]));
    L6MUX21 i12287 (.D0(n15947), .D1(n15948), .SD(raddr13_ff), .Z(Sprite_readData[5]));
    L6MUX21 i12302 (.D0(n15962), .D1(n15963), .SD(raddr13_ff), .Z(Sprite_readData[6]));
    L6MUX21 i12317 (.D0(n15977), .D1(n15978), .SD(raddr13_ff), .Z(Sprite_readData[7]));
    LUT4 i12215_3_lut (.A(mdout1_4_1), .B(mdout1_5_1), .C(raddr10_ff), 
         .Z(n15877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12215_3_lut.init = 16'hcaca;
    L6MUX21 i12332 (.D0(n15992), .D1(n15993), .SD(raddr13_ff), .Z(Sprite_readData[8]));
    L6MUX21 i12212 (.D0(n15872), .D1(n15873), .SD(raddr13_ff), .Z(Sprite_readData[0]));
    L6MUX21 i12227 (.D0(n15887), .D1(n15888), .SD(raddr13_ff), .Z(Sprite_readData[1]));
    L6MUX21 i12241 (.D0(n15900), .D1(n15901), .SD(raddr12_ff), .Z(n15903));
    L6MUX21 i12255 (.D0(n15913), .D1(n15914), .SD(raddr12_ff), .Z(n15917));
    L6MUX21 i12256 (.D0(n15915), .D1(n15916), .SD(raddr12_ff), .Z(n15918));
    L6MUX21 i12270 (.D0(n15928), .D1(n15929), .SD(raddr12_ff), .Z(n15932));
    L6MUX21 i12271 (.D0(n15930), .D1(n15931), .SD(raddr12_ff), .Z(n15933));
    L6MUX21 i12285 (.D0(n15943), .D1(n15944), .SD(raddr12_ff), .Z(n15947));
    L6MUX21 i12286 (.D0(n15945), .D1(n15946), .SD(raddr12_ff), .Z(n15948));
    L6MUX21 i12300 (.D0(n15958), .D1(n15959), .SD(raddr12_ff), .Z(n15962));
    L6MUX21 i12301 (.D0(n15960), .D1(n15961), .SD(raddr12_ff), .Z(n15963));
    L6MUX21 i12315 (.D0(n15973), .D1(n15974), .SD(raddr12_ff), .Z(n15977));
    L6MUX21 i12316 (.D0(n15975), .D1(n15976), .SD(raddr12_ff), .Z(n15978));
    L6MUX21 i12330 (.D0(n15988), .D1(n15989), .SD(raddr12_ff), .Z(n15992));
    L6MUX21 i12331 (.D0(n15990), .D1(n15991), .SD(raddr12_ff), .Z(n15993));
    LUT4 i12201_3_lut (.A(mdout1_6_0), .B(mdout1_7_0), .C(raddr10_ff), 
         .Z(n15863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12201_3_lut.init = 16'hcaca;
    LUT4 i12214_3_lut (.A(mdout1_2_1), .B(mdout1_3_1), .C(raddr10_ff), 
         .Z(n15876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12214_3_lut.init = 16'hcaca;
    L6MUX21 i12210 (.D0(n15868), .D1(n15869), .SD(raddr12_ff), .Z(n15872));
    PFUMX i12238 (.BLUT(n15894), .ALUT(n15895), .C0(raddr11_ff), .Z(n15900));
    L6MUX21 i12211 (.D0(n15870), .D1(n15871), .SD(raddr12_ff), .Z(n15873));
    L6MUX21 i12225 (.D0(n15883), .D1(n15884), .SD(raddr12_ff), .Z(n15887));
    L6MUX21 i12226 (.D0(n15885), .D1(n15886), .SD(raddr12_ff), .Z(n15888));
    L6MUX21 i12240 (.D0(n15898), .D1(n15899), .SD(raddr12_ff), .Z(n15902));
    PFUMX i12251 (.BLUT(n15905), .ALUT(n15906), .C0(raddr11_ff), .Z(n15913));
    PFUMX i12252 (.BLUT(n15907), .ALUT(n15908), .C0(raddr11_ff), .Z(n15914));
    PFUMX i12253 (.BLUT(n15909), .ALUT(n15910), .C0(raddr11_ff), .Z(n15915));
    PFUMX i12254 (.BLUT(n15911), .ALUT(n15912), .C0(raddr11_ff), .Z(n15916));
    PFUMX i12266 (.BLUT(n15920), .ALUT(n15921), .C0(raddr11_ff), .Z(n15928));
    PFUMX i12267 (.BLUT(n15922), .ALUT(n15923), .C0(raddr11_ff), .Z(n15929));
    PFUMX i12268 (.BLUT(n15924), .ALUT(n15925), .C0(raddr11_ff), .Z(n15930));
    PFUMX i12269 (.BLUT(n15926), .ALUT(n15927), .C0(raddr11_ff), .Z(n15931));
    LUT4 i12213_3_lut (.A(mdout1_0_1), .B(mdout1_1_1), .C(raddr10_ff), 
         .Z(n15875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12213_3_lut.init = 16'hcaca;
    PFUMX i12281 (.BLUT(n15935), .ALUT(n15936), .C0(raddr11_ff), .Z(n15943));
    PFUMX i12282 (.BLUT(n15937), .ALUT(n15938), .C0(raddr11_ff), .Z(n15944));
    PFUMX i12283 (.BLUT(n15939), .ALUT(n15940), .C0(raddr11_ff), .Z(n15945));
    LUT4 i12199_3_lut (.A(mdout1_2_0), .B(mdout1_3_0), .C(raddr10_ff), 
         .Z(n15861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12199_3_lut.init = 16'hcaca;
    LUT4 i12229_3_lut (.A(mdout1_2_2), .B(mdout1_3_2), .C(raddr10_ff), 
         .Z(n15891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12229_3_lut.init = 16'hcaca;
    PFUMX i12284 (.BLUT(n15941), .ALUT(n15942), .C0(raddr11_ff), .Z(n15946));
    PFUMX i12296 (.BLUT(n15950), .ALUT(n15951), .C0(raddr11_ff), .Z(n15958));
    PFUMX i12297 (.BLUT(n15952), .ALUT(n15953), .C0(raddr11_ff), .Z(n15959));
    PFUMX i12298 (.BLUT(n15954), .ALUT(n15955), .C0(raddr11_ff), .Z(n15960));
    PFUMX i12299 (.BLUT(n15956), .ALUT(n15957), .C0(raddr11_ff), .Z(n15961));
    PFUMX i12311 (.BLUT(n15965), .ALUT(n15966), .C0(raddr11_ff), .Z(n15973));
    PFUMX i12312 (.BLUT(n15967), .ALUT(n15968), .C0(raddr11_ff), .Z(n15974));
    PFUMX i12313 (.BLUT(n15969), .ALUT(n15970), .C0(raddr11_ff), .Z(n15975));
    PFUMX i12314 (.BLUT(n15971), .ALUT(n15972), .C0(raddr11_ff), .Z(n15976));
    PFUMX i12326 (.BLUT(n15980), .ALUT(n15981), .C0(raddr11_ff), .Z(n15988));
    PFUMX i12327 (.BLUT(n15982), .ALUT(n15983), .C0(raddr11_ff), .Z(n15989));
    PFUMX i12328 (.BLUT(n15984), .ALUT(n15985), .C0(raddr11_ff), .Z(n15990));
    PFUMX i12329 (.BLUT(n15986), .ALUT(n15987), .C0(raddr11_ff), .Z(n15991));
    PFUMX i12239 (.BLUT(n15896), .ALUT(n15897), .C0(raddr11_ff), .Z(n15901));
    LUT4 i12198_3_lut (.A(mdout1_0_0), .B(mdout1_1_0), .C(raddr10_ff), 
         .Z(n15860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12198_3_lut.init = 16'hcaca;
    LUT4 i12228_3_lut (.A(mdout1_0_2), .B(mdout1_1_2), .C(raddr10_ff), 
         .Z(n15890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12228_3_lut.init = 16'hcaca;
    PFUMX i12223 (.BLUT(n15879), .ALUT(n15880), .C0(raddr11_ff), .Z(n15885));
    LUT4 i12220_3_lut (.A(mdout1_14_1), .B(mdout1_15_1), .C(raddr10_ff), 
         .Z(n15882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12220_3_lut.init = 16'hcaca;
    LUT4 i12205_3_lut (.A(mdout1_14_0), .B(mdout1_15_0), .C(raddr10_ff), 
         .Z(n15867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12205_3_lut.init = 16'hcaca;
    LUT4 i12204_3_lut (.A(mdout1_12_0), .B(mdout1_13_0), .C(raddr10_ff), 
         .Z(n15866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12204_3_lut.init = 16'hcaca;
    LUT4 i12203_3_lut (.A(mdout1_10_0), .B(mdout1_11_0), .C(raddr10_ff), 
         .Z(n15865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12203_3_lut.init = 16'hcaca;
    LUT4 i12202_3_lut (.A(mdout1_8_0), .B(mdout1_9_0), .C(raddr10_ff), 
         .Z(n15864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12202_3_lut.init = 16'hcaca;
    LUT4 i12219_3_lut (.A(mdout1_12_1), .B(mdout1_13_1), .C(raddr10_ff), 
         .Z(n15881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(634[8:17])
    defparam i12219_3_lut.init = 16'hcaca;
    PFUMX i12224 (.BLUT(n15881), .ALUT(n15882), .C0(raddr11_ff), .Z(n15886));
    
endmodule
//
// Verilog Description of module LUT_RAM
//

module LUT_RAM (\BUS_data[8] , \BUS_data[7] , \BUS_data[6] , \BUS_data[5] , 
            \BUS_data[4] , \BUS_data[3] , \BUS_data[2] , \BUS_data[1] , 
            \BUS_data[0] , GND_net, \BUS_addr[10] , n17325, n17337, 
            n17334, n17321, n17331, n17332, n17333, n17339, Sprite_readData, 
            SpriteLut_writeClk, SpriteLut_readClk, VCC_net, RED_WE, 
            RED_WRITE, RED_READ) /* synthesis NGD_DRC_MASK=1 */ ;
    input \BUS_data[8] ;
    input \BUS_data[7] ;
    input \BUS_data[6] ;
    input \BUS_data[5] ;
    input \BUS_data[4] ;
    input \BUS_data[3] ;
    input \BUS_data[2] ;
    input \BUS_data[1] ;
    input \BUS_data[0] ;
    input GND_net;
    input \BUS_addr[10] ;
    input n17325;
    input n17337;
    input n17334;
    input n17321;
    input n17331;
    input n17332;
    input n17333;
    input n17339;
    input [8:0]Sprite_readData;
    input SpriteLut_writeClk;
    input SpriteLut_readClk;
    input VCC_net;
    input RED_WE;
    output [8:0]RED_WRITE;
    output [8:0]RED_READ;
    
    wire SpriteLut_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(202[9:27])
    wire SpriteLut_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(203[9:26])
    
    DP8KC LUT_RAM_0_0_0 (.DIA0(\BUS_data[0] ), .DIA1(\BUS_data[1] ), .DIA2(\BUS_data[2] ), 
          .DIA3(\BUS_data[3] ), .DIA4(\BUS_data[4] ), .DIA5(\BUS_data[5] ), 
          .DIA6(\BUS_data[6] ), .DIA7(\BUS_data[7] ), .DIA8(\BUS_data[8] ), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(n17339), 
          .ADA4(n17333), .ADA5(n17332), .ADA6(n17331), .ADA7(n17321), 
          .ADA8(n17334), .ADA9(n17337), .ADA10(n17325), .ADA11(\BUS_addr[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(SpriteLut_writeClk), 
          .WEA(RED_WE), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(Sprite_readData[0]), .ADB4(Sprite_readData[1]), 
          .ADB5(Sprite_readData[2]), .ADB6(Sprite_readData[3]), .ADB7(Sprite_readData[4]), 
          .ADB8(Sprite_readData[5]), .ADB9(Sprite_readData[6]), .ADB10(Sprite_readData[7]), 
          .ADB11(Sprite_readData[8]), .ADB12(GND_net), .CEB(VCC_net), 
          .OCEB(VCC_net), .CLKB(SpriteLut_readClk), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOA0(RED_WRITE[0]), 
          .DOA1(RED_WRITE[1]), .DOA2(RED_WRITE[2]), .DOA3(RED_WRITE[3]), 
          .DOA4(RED_WRITE[4]), .DOA5(RED_WRITE[5]), .DOA6(RED_WRITE[6]), 
          .DOA7(RED_WRITE[7]), .DOA8(RED_WRITE[8]), .DOB0(RED_READ[0]), 
          .DOB1(RED_READ[1]), .DOB2(RED_READ[2]), .DOB3(RED_READ[3]), 
          .DOB4(RED_READ[4]), .DOB5(RED_READ[5]), .DOB6(RED_READ[6]), 
          .DOB7(RED_READ[7]), .DOB8(RED_READ[8])) /* synthesis MEM_LPC_FILE="LUT_RAM.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=11, LSE_RCOL=18, LSE_LLINE=651, LSE_RLINE=651 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(651[11:18])
    defparam LUT_RAM_0_0_0.DATA_WIDTH_A = 9;
    defparam LUT_RAM_0_0_0.DATA_WIDTH_B = 9;
    defparam LUT_RAM_0_0_0.REGMODE_A = "NOREG";
    defparam LUT_RAM_0_0_0.REGMODE_B = "NOREG";
    defparam LUT_RAM_0_0_0.CSDECODE_A = "0b000";
    defparam LUT_RAM_0_0_0.CSDECODE_B = "0b000";
    defparam LUT_RAM_0_0_0.WRITEMODE_A = "NORMAL";
    defparam LUT_RAM_0_0_0.WRITEMODE_B = "NORMAL";
    defparam LUT_RAM_0_0_0.GSR = "ENABLED";
    defparam LUT_RAM_0_0_0.RESETMODE = "ASYNC";
    defparam LUT_RAM_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam LUT_RAM_0_0_0.INIT_DATA = "STATIC";
    defparam LUT_RAM_0_0_0.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    
endmodule
//
// Verilog Description of module LUT_RAM_U0
//

module LUT_RAM_U0 (\BUS_data[8] , \BUS_data[7] , \BUS_data[6] , \BUS_data[5] , 
            \BUS_data[4] , \BUS_data[3] , \BUS_data[2] , \BUS_data[1] , 
            \BUS_data[0] , GND_net, \BUS_addr[10] , n17325, n17337, 
            n17334, n17321, n17331, n17332, n17333, n17339, Sprite_readData, 
            SpriteLut_writeClk, SpriteLut_readClk, VCC_net, GREEN_WE, 
            GREEN_WRITE, GREEN_READ) /* synthesis NGD_DRC_MASK=1 */ ;
    input \BUS_data[8] ;
    input \BUS_data[7] ;
    input \BUS_data[6] ;
    input \BUS_data[5] ;
    input \BUS_data[4] ;
    input \BUS_data[3] ;
    input \BUS_data[2] ;
    input \BUS_data[1] ;
    input \BUS_data[0] ;
    input GND_net;
    input \BUS_addr[10] ;
    input n17325;
    input n17337;
    input n17334;
    input n17321;
    input n17331;
    input n17332;
    input n17333;
    input n17339;
    input [8:0]Sprite_readData;
    input SpriteLut_writeClk;
    input SpriteLut_readClk;
    input VCC_net;
    input GREEN_WE;
    output [8:0]GREEN_WRITE;
    output [8:0]GREEN_READ;
    
    wire SpriteLut_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(202[9:27])
    wire SpriteLut_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(203[9:26])
    
    DP8KC LUT_RAM_0_0_0 (.DIA0(\BUS_data[0] ), .DIA1(\BUS_data[1] ), .DIA2(\BUS_data[2] ), 
          .DIA3(\BUS_data[3] ), .DIA4(\BUS_data[4] ), .DIA5(\BUS_data[5] ), 
          .DIA6(\BUS_data[6] ), .DIA7(\BUS_data[7] ), .DIA8(\BUS_data[8] ), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(n17339), 
          .ADA4(n17333), .ADA5(n17332), .ADA6(n17331), .ADA7(n17321), 
          .ADA8(n17334), .ADA9(n17337), .ADA10(n17325), .ADA11(\BUS_addr[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(SpriteLut_writeClk), 
          .WEA(GREEN_WE), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(Sprite_readData[0]), .ADB4(Sprite_readData[1]), 
          .ADB5(Sprite_readData[2]), .ADB6(Sprite_readData[3]), .ADB7(Sprite_readData[4]), 
          .ADB8(Sprite_readData[5]), .ADB9(Sprite_readData[6]), .ADB10(Sprite_readData[7]), 
          .ADB11(Sprite_readData[8]), .ADB12(GND_net), .CEB(VCC_net), 
          .OCEB(VCC_net), .CLKB(SpriteLut_readClk), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOA0(GREEN_WRITE[0]), 
          .DOA1(GREEN_WRITE[1]), .DOA2(GREEN_WRITE[2]), .DOA3(GREEN_WRITE[3]), 
          .DOA4(GREEN_WRITE[4]), .DOA5(GREEN_WRITE[5]), .DOA6(GREEN_WRITE[6]), 
          .DOA7(GREEN_WRITE[7]), .DOA8(GREEN_WRITE[8]), .DOB0(GREEN_READ[0]), 
          .DOB1(GREEN_READ[1]), .DOB2(GREEN_READ[2]), .DOB3(GREEN_READ[3]), 
          .DOB4(GREEN_READ[4]), .DOB5(GREEN_READ[5]), .DOB6(GREEN_READ[6]), 
          .DOB7(GREEN_READ[7]), .DOB8(GREEN_READ[8])) /* synthesis MEM_LPC_FILE="LUT_RAM.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=12, LSE_RCOL=19, LSE_LLINE=669, LSE_RLINE=669 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(669[12:19])
    defparam LUT_RAM_0_0_0.DATA_WIDTH_A = 9;
    defparam LUT_RAM_0_0_0.DATA_WIDTH_B = 9;
    defparam LUT_RAM_0_0_0.REGMODE_A = "NOREG";
    defparam LUT_RAM_0_0_0.REGMODE_B = "NOREG";
    defparam LUT_RAM_0_0_0.CSDECODE_A = "0b000";
    defparam LUT_RAM_0_0_0.CSDECODE_B = "0b000";
    defparam LUT_RAM_0_0_0.WRITEMODE_A = "NORMAL";
    defparam LUT_RAM_0_0_0.WRITEMODE_B = "NORMAL";
    defparam LUT_RAM_0_0_0.GSR = "ENABLED";
    defparam LUT_RAM_0_0_0.RESETMODE = "ASYNC";
    defparam LUT_RAM_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam LUT_RAM_0_0_0.INIT_DATA = "STATIC";
    defparam LUT_RAM_0_0_0.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    
endmodule
//
// Verilog Description of module GammaRam
//

module GammaRam (\BUS_data[9] , GND_net, GR_WR_ADDR, currValue, GR_WR_CLK, 
            LOGIC_CLOCK_N_57, VCC_net, n17387, GR_WR_DOUT, GR_RE_DOUT, 
            \BUS_data[8] , \BUS_data[7] , \BUS_data[6] , \BUS_data[5] , 
            \BUS_data[4] , \BUS_data[3] , \BUS_data[2] , \BUS_data[1] , 
            \BUS_data[0] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input \BUS_data[9] ;
    input GND_net;
    input [7:0]GR_WR_ADDR;
    input [7:0]currValue;
    input GR_WR_CLK;
    input LOGIC_CLOCK_N_57;
    input VCC_net;
    input n17387;
    output [9:0]GR_WR_DOUT;
    output [9:0]GR_RE_DOUT;
    input \BUS_data[8] ;
    input \BUS_data[7] ;
    input \BUS_data[6] ;
    input \BUS_data[5] ;
    input \BUS_data[4] ;
    input \BUS_data[3] ;
    input \BUS_data[2] ;
    input \BUS_data[1] ;
    input \BUS_data[0] ;
    
    wire GR_WR_CLK /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(162[9:18])
    wire LOGIC_CLOCK_N_57 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    
    DP8KC GammaRam_0_1_0 (.DIA0(\BUS_data[9] ), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(GR_WR_ADDR[0]), .ADA4(GR_WR_ADDR[1]), 
          .ADA5(GR_WR_ADDR[2]), .ADA6(GR_WR_ADDR[3]), .ADA7(GR_WR_ADDR[4]), 
          .ADA8(GR_WR_ADDR[5]), .ADA9(GR_WR_ADDR[6]), .ADA10(GR_WR_ADDR[7]), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(GR_WR_CLK), .WEA(n17387), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(currValue[0]), .ADB4(currValue[1]), 
          .ADB5(currValue[2]), .ADB6(currValue[3]), .ADB7(currValue[4]), 
          .ADB8(currValue[5]), .ADB9(currValue[6]), .ADB10(currValue[7]), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(LOGIC_CLOCK_N_57), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(GR_WR_DOUT[9]), .DOB0(GR_RE_DOUT[9])) /* synthesis MEM_LPC_FILE="GammaRam.lpc", MEM_INIT_FILE="gammadefault.mem", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=16, LSE_LLINE=616, LSE_RLINE=616 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(616[8:16])
    defparam GammaRam_0_1_0.DATA_WIDTH_A = 9;
    defparam GammaRam_0_1_0.DATA_WIDTH_B = 9;
    defparam GammaRam_0_1_0.REGMODE_A = "NOREG";
    defparam GammaRam_0_1_0.REGMODE_B = "NOREG";
    defparam GammaRam_0_1_0.CSDECODE_A = "0b000";
    defparam GammaRam_0_1_0.CSDECODE_B = "0b000";
    defparam GammaRam_0_1_0.WRITEMODE_A = "NORMAL";
    defparam GammaRam_0_1_0.WRITEMODE_B = "NORMAL";
    defparam GammaRam_0_1_0.GSR = "ENABLED";
    defparam GammaRam_0_1_0.RESETMODE = "ASYNC";
    defparam GammaRam_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam GammaRam_0_1_0.INIT_DATA = "STATIC";
    defparam GammaRam_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_04 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_05 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_06 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_07 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC GammaRam_0_0_1 (.DIA0(\BUS_data[0] ), .DIA1(\BUS_data[1] ), .DIA2(\BUS_data[2] ), 
          .DIA3(\BUS_data[3] ), .DIA4(\BUS_data[4] ), .DIA5(\BUS_data[5] ), 
          .DIA6(\BUS_data[6] ), .DIA7(\BUS_data[7] ), .DIA8(\BUS_data[8] ), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(GR_WR_ADDR[0]), 
          .ADA4(GR_WR_ADDR[1]), .ADA5(GR_WR_ADDR[2]), .ADA6(GR_WR_ADDR[3]), 
          .ADA7(GR_WR_ADDR[4]), .ADA8(GR_WR_ADDR[5]), .ADA9(GR_WR_ADDR[6]), 
          .ADA10(GR_WR_ADDR[7]), .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), 
          .OCEA(VCC_net), .CLKA(GR_WR_CLK), .WEA(n17387), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(VCC_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(currValue[0]), 
          .ADB4(currValue[1]), .ADB5(currValue[2]), .ADB6(currValue[3]), 
          .ADB7(currValue[4]), .ADB8(currValue[5]), .ADB9(currValue[6]), 
          .ADB10(currValue[7]), .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), 
          .OCEB(VCC_net), .CLKB(LOGIC_CLOCK_N_57), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOA0(GR_WR_DOUT[0]), 
          .DOA1(GR_WR_DOUT[1]), .DOA2(GR_WR_DOUT[2]), .DOA3(GR_WR_DOUT[3]), 
          .DOA4(GR_WR_DOUT[4]), .DOA5(GR_WR_DOUT[5]), .DOA6(GR_WR_DOUT[6]), 
          .DOA7(GR_WR_DOUT[7]), .DOA8(GR_WR_DOUT[8]), .DOB0(GR_RE_DOUT[0]), 
          .DOB1(GR_RE_DOUT[1]), .DOB2(GR_RE_DOUT[2]), .DOB3(GR_RE_DOUT[3]), 
          .DOB4(GR_RE_DOUT[4]), .DOB5(GR_RE_DOUT[5]), .DOB6(GR_RE_DOUT[6]), 
          .DOB7(GR_RE_DOUT[7]), .DOB8(GR_RE_DOUT[8])) /* synthesis MEM_LPC_FILE="GammaRam.lpc", MEM_INIT_FILE="gammadefault.mem", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=16, LSE_LLINE=616, LSE_RLINE=616 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(616[8:16])
    defparam GammaRam_0_0_1.DATA_WIDTH_A = 9;
    defparam GammaRam_0_0_1.DATA_WIDTH_B = 9;
    defparam GammaRam_0_0_1.REGMODE_A = "NOREG";
    defparam GammaRam_0_0_1.REGMODE_B = "NOREG";
    defparam GammaRam_0_0_1.CSDECODE_A = "0b000";
    defparam GammaRam_0_0_1.CSDECODE_B = "0b000";
    defparam GammaRam_0_0_1.WRITEMODE_A = "NORMAL";
    defparam GammaRam_0_0_1.WRITEMODE_B = "NORMAL";
    defparam GammaRam_0_0_1.GSR = "ENABLED";
    defparam GammaRam_0_0_1.RESETMODE = "ASYNC";
    defparam GammaRam_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam GammaRam_0_0_1.INIT_DATA = "STATIC";
    defparam GammaRam_0_0_1.INITVAL_00 = "0x0F8780E8700D8680C8600B8580A85009848088400783806830058280482003818028100180800800";
    defparam GammaRam_0_0_1.INITVAL_01 = "0x1F8F81E8F01D8E81C8E01B8D81A8D0198C8188C0178B8168B0158A8148A013898128901188810880";
    defparam GammaRam_0_0_1.INITVAL_02 = "0x2F9782E9702D9682C9602B9582A95029948289402793826930259282492023918229102190820900";
    defparam GammaRam_0_0_1.INITVAL_03 = "0x3F9F83E9F03D9E83C9E03B9D83A9D0399C8389C0379B8369B0359A8349A033998329903198830980";
    defparam GammaRam_0_0_1.INITVAL_04 = "0x0F8780E8700D8680C8600B8580A85009848088400783806830058280482003818028100180800800";
    defparam GammaRam_0_0_1.INITVAL_05 = "0x1F8F81E8F01D8E81C8E01B8D81A8D0198C8188C0178B8168B0158A8148A013898128901188810880";
    defparam GammaRam_0_0_1.INITVAL_06 = "0x2F9782E9702D9682C9602B9582A95029948289402793826930259282492023918229102190820900";
    defparam GammaRam_0_0_1.INITVAL_07 = "0x3F9F83E9F03D9E83C9E03B9D83A9D0399C8389C0379B8369B0359A8349A033998329903198830980";
    defparam GammaRam_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module LUT_RAM_U1
//

module LUT_RAM_U1 (\BUS_data[8] , \BUS_data[7] , \BUS_data[6] , \BUS_data[5] , 
            \BUS_data[4] , \BUS_data[3] , \BUS_data[2] , \BUS_data[1] , 
            \BUS_data[0] , GND_net, \BUS_addr[10] , n17325, n17337, 
            n17334, n17321, n17331, n17332, n17333, n17339, Sprite_readData, 
            SpriteLut_writeClk, SpriteLut_readClk, VCC_net, BLUE_WE, 
            BLUE_WRITE, BLUE_READ) /* synthesis NGD_DRC_MASK=1 */ ;
    input \BUS_data[8] ;
    input \BUS_data[7] ;
    input \BUS_data[6] ;
    input \BUS_data[5] ;
    input \BUS_data[4] ;
    input \BUS_data[3] ;
    input \BUS_data[2] ;
    input \BUS_data[1] ;
    input \BUS_data[0] ;
    input GND_net;
    input \BUS_addr[10] ;
    input n17325;
    input n17337;
    input n17334;
    input n17321;
    input n17331;
    input n17332;
    input n17333;
    input n17339;
    input [8:0]Sprite_readData;
    input SpriteLut_writeClk;
    input SpriteLut_readClk;
    input VCC_net;
    input BLUE_WE;
    output [8:0]BLUE_WRITE;
    output [8:0]BLUE_READ;
    
    wire SpriteLut_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(202[9:27])
    wire SpriteLut_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(203[9:26])
    
    DP8KC LUT_RAM_0_0_0 (.DIA0(\BUS_data[0] ), .DIA1(\BUS_data[1] ), .DIA2(\BUS_data[2] ), 
          .DIA3(\BUS_data[3] ), .DIA4(\BUS_data[4] ), .DIA5(\BUS_data[5] ), 
          .DIA6(\BUS_data[6] ), .DIA7(\BUS_data[7] ), .DIA8(\BUS_data[8] ), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(n17339), 
          .ADA4(n17333), .ADA5(n17332), .ADA6(n17331), .ADA7(n17321), 
          .ADA8(n17334), .ADA9(n17337), .ADA10(n17325), .ADA11(\BUS_addr[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(SpriteLut_writeClk), 
          .WEA(BLUE_WE), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(Sprite_readData[0]), .ADB4(Sprite_readData[1]), 
          .ADB5(Sprite_readData[2]), .ADB6(Sprite_readData[3]), .ADB7(Sprite_readData[4]), 
          .ADB8(Sprite_readData[5]), .ADB9(Sprite_readData[6]), .ADB10(Sprite_readData[7]), 
          .ADB11(Sprite_readData[8]), .ADB12(GND_net), .CEB(VCC_net), 
          .OCEB(VCC_net), .CLKB(SpriteLut_readClk), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOA0(BLUE_WRITE[0]), 
          .DOA1(BLUE_WRITE[1]), .DOA2(BLUE_WRITE[2]), .DOA3(BLUE_WRITE[3]), 
          .DOA4(BLUE_WRITE[4]), .DOA5(BLUE_WRITE[5]), .DOA6(BLUE_WRITE[6]), 
          .DOA7(BLUE_WRITE[7]), .DOA8(BLUE_WRITE[8]), .DOB0(BLUE_READ[0]), 
          .DOB1(BLUE_READ[1]), .DOB2(BLUE_READ[2]), .DOB3(BLUE_READ[3]), 
          .DOB4(BLUE_READ[4]), .DOB5(BLUE_READ[5]), .DOB6(BLUE_READ[6]), 
          .DOB7(BLUE_READ[7]), .DOB8(BLUE_READ[8])) /* synthesis MEM_LPC_FILE="LUT_RAM.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=11, LSE_RCOL=18, LSE_LLINE=687, LSE_RLINE=687 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(687[11:18])
    defparam LUT_RAM_0_0_0.DATA_WIDTH_A = 9;
    defparam LUT_RAM_0_0_0.DATA_WIDTH_B = 9;
    defparam LUT_RAM_0_0_0.REGMODE_A = "NOREG";
    defparam LUT_RAM_0_0_0.REGMODE_B = "NOREG";
    defparam LUT_RAM_0_0_0.CSDECODE_A = "0b000";
    defparam LUT_RAM_0_0_0.CSDECODE_B = "0b000";
    defparam LUT_RAM_0_0_0.WRITEMODE_A = "NORMAL";
    defparam LUT_RAM_0_0_0.WRITEMODE_B = "NORMAL";
    defparam LUT_RAM_0_0_0.GSR = "ENABLED";
    defparam LUT_RAM_0_0_0.RESETMODE = "ASYNC";
    defparam LUT_RAM_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam LUT_RAM_0_0_0.INIT_DATA = "STATIC";
    defparam LUT_RAM_0_0_0.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    
endmodule
//
// Verilog Description of module LUT_RAM_U2
//

module LUT_RAM_U2 (\BUS_data[8] , \BUS_data[7] , \BUS_data[6] , \BUS_data[5] , 
            \BUS_data[4] , \BUS_data[3] , \BUS_data[2] , \BUS_data[1] , 
            \BUS_data[0] , GND_net, \BUS_addr[10] , n17325, n17337, 
            n17334, n17321, n17331, n17332, n17333, n17339, Sprite_readData, 
            SpriteLut_writeClk, SpriteLut_readClk, VCC_net, ALPHA_WE, 
            ALPHA_WRITE, ALPHA_READ) /* synthesis NGD_DRC_MASK=1 */ ;
    input \BUS_data[8] ;
    input \BUS_data[7] ;
    input \BUS_data[6] ;
    input \BUS_data[5] ;
    input \BUS_data[4] ;
    input \BUS_data[3] ;
    input \BUS_data[2] ;
    input \BUS_data[1] ;
    input \BUS_data[0] ;
    input GND_net;
    input \BUS_addr[10] ;
    input n17325;
    input n17337;
    input n17334;
    input n17321;
    input n17331;
    input n17332;
    input n17333;
    input n17339;
    input [8:0]Sprite_readData;
    input SpriteLut_writeClk;
    input SpriteLut_readClk;
    input VCC_net;
    input ALPHA_WE;
    output [8:0]ALPHA_WRITE;
    output [8:0]ALPHA_READ;
    
    wire SpriteLut_writeClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(202[9:27])
    wire SpriteLut_readClk /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(203[9:26])
    
    DP8KC LUT_RAM_0_0_0 (.DIA0(\BUS_data[0] ), .DIA1(\BUS_data[1] ), .DIA2(\BUS_data[2] ), 
          .DIA3(\BUS_data[3] ), .DIA4(\BUS_data[4] ), .DIA5(\BUS_data[5] ), 
          .DIA6(\BUS_data[6] ), .DIA7(\BUS_data[7] ), .DIA8(\BUS_data[8] ), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(n17339), 
          .ADA4(n17333), .ADA5(n17332), .ADA6(n17331), .ADA7(n17321), 
          .ADA8(n17334), .ADA9(n17337), .ADA10(n17325), .ADA11(\BUS_addr[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(SpriteLut_writeClk), 
          .WEA(ALPHA_WE), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(Sprite_readData[0]), .ADB4(Sprite_readData[1]), 
          .ADB5(Sprite_readData[2]), .ADB6(Sprite_readData[3]), .ADB7(Sprite_readData[4]), 
          .ADB8(Sprite_readData[5]), .ADB9(Sprite_readData[6]), .ADB10(Sprite_readData[7]), 
          .ADB11(Sprite_readData[8]), .ADB12(GND_net), .CEB(VCC_net), 
          .OCEB(VCC_net), .CLKB(SpriteLut_readClk), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOA0(ALPHA_WRITE[0]), 
          .DOA1(ALPHA_WRITE[1]), .DOA2(ALPHA_WRITE[2]), .DOA3(ALPHA_WRITE[3]), 
          .DOA4(ALPHA_WRITE[4]), .DOA5(ALPHA_WRITE[5]), .DOA6(ALPHA_WRITE[6]), 
          .DOA7(ALPHA_WRITE[7]), .DOA8(ALPHA_WRITE[8]), .DOB0(ALPHA_READ[0]), 
          .DOB1(ALPHA_READ[1]), .DOB2(ALPHA_READ[2]), .DOB3(ALPHA_READ[3]), 
          .DOB4(ALPHA_READ[4]), .DOB5(ALPHA_READ[5]), .DOB6(ALPHA_READ[6]), 
          .DOB7(ALPHA_READ[7]), .DOB8(ALPHA_READ[8])) /* synthesis MEM_LPC_FILE="LUT_RAM.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=12, LSE_RCOL=19, LSE_LLINE=705, LSE_RLINE=705 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(705[12:19])
    defparam LUT_RAM_0_0_0.DATA_WIDTH_A = 9;
    defparam LUT_RAM_0_0_0.DATA_WIDTH_B = 9;
    defparam LUT_RAM_0_0_0.REGMODE_A = "NOREG";
    defparam LUT_RAM_0_0_0.REGMODE_B = "NOREG";
    defparam LUT_RAM_0_0_0.CSDECODE_A = "0b000";
    defparam LUT_RAM_0_0_0.CSDECODE_B = "0b000";
    defparam LUT_RAM_0_0_0.WRITEMODE_A = "NORMAL";
    defparam LUT_RAM_0_0_0.WRITEMODE_B = "NORMAL";
    defparam LUT_RAM_0_0_0.GSR = "ENABLED";
    defparam LUT_RAM_0_0_0.RESETMODE = "ASYNC";
    defparam LUT_RAM_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam LUT_RAM_0_0_0.INIT_DATA = "STATIC";
    defparam LUT_RAM_0_0_0.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam LUT_RAM_0_0_0.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    
endmodule
//
// Verilog Description of module PIC
//

module PIC (PIC_DATA_IN_out_7, \BUS_currGrantID[1] , \BUS_currGrantID[0] , 
            \BUS_ADDR_INTERNAL[11] , n18273, \BUS_ADDR_INTERNAL[12] , 
            n18272, GND_net, writeData, LOGIC_CLOCK, PIC_DATA_IN_out_15, 
            PIC_DATA_IN_out_14, PIC_DATA_IN_out_13, PIC_DATA_IN_out_12, 
            PIC_DATA_IN_out_11, \BUS_ADDR_INTERNAL[9] , n18268, \BUS_ADDR_INTERNAL[10] , 
            n18269, \BUS_ADDR_INTERNAL[8] , n18267, OUT_ENABLE, n9950, 
            \PIC_data[0] , \writeData[10] , PIC_DATA_IN_out_10, \writeData[9] , 
            PIC_DATA_IN_out_9, \writeData[8] , PIC_DATA_IN_out_8, n17298, 
            n17337, n17325, n15534, state, n17270, PIC_WE_IN_c, 
            \BUS_data[0] , \BUS_ADDR_INTERNAL[0] , PIC_ADDR_IN_c_0, \BUS_ADDR_INTERNAL[1] , 
            \BUS_ADDR_INTERNAL[1]_adj_1 , n17384, \BUS_req[2] , \BUS_ADDR_INTERNAL[18] , 
            n2642, LOGIC_CLOCK_enable_52, n2504, n17279, PIC_DATA_IN_out_0, 
            WRITE_DONE, n18280, PIC_ADDR_IN_c_1, PIC_ADDR_IN_c_2, PIC_ADDR_IN_c_3, 
            PIC_ADDR_IN_c_4, PIC_ADDR_IN_c_5, PIC_ADDR_IN_c_6, PIC_ADDR_IN_c_7, 
            PIC_ADDR_IN_c_8, PIC_ADDR_IN_c_9, PIC_ADDR_IN_c_10, PIC_ADDR_IN_c_11, 
            PIC_ADDR_IN_c_12, PIC_ADDR_IN_c_13, PIC_ADDR_IN_c_14, PIC_ADDR_IN_c_15, 
            PIC_ADDR_IN_c_16, PIC_ADDR_IN_c_17, PIC_ADDR_IN_c_18, n14, 
            n17434, BUS_DIRECTION_INTERNAL, n18260, n16456, n17276, 
            LOGIC_CLOCK_N_57_enable_3, n17457, n17278, n15571, PIC_OE_c, 
            n15469, PIC_READY_c, SpriteRead_yInSprite, \currSprite_size[6] , 
            \currSprite_size[4] , \currSprite_size[2] , n17394, \Sprite_readAddr_13__N_752[0] , 
            \Sprite_readAddr_13__N_752[2] , \Sprite_readAddr_13__N_752[3] , 
            \Sprite_readAddr_13__N_752[4] , \Sprite_readAddr_13__N_752[6] , 
            \Sprite_readAddr_13__N_752[5] , \Sprite_readAddr_13__N_752[8] , 
            \Sprite_readAddr_13__N_752[7] , \Sprite_readAddr_13__N_752[10] , 
            \Sprite_readAddr_13__N_752[9] , \Sprite_readAddr_13__N_752[12] , 
            \Sprite_readAddr_13__N_752[11] , \Sprite_readAddr_13__N_752[13] , 
            \currSprite_size[1] , \Sprite_readAddr_13__N_752[1] , \currSprite_size[3] , 
            \currSprite_size[5] , \currSprite_size[7] , \BUS_data[1] , 
            \BUS_data[2] , \BUS_data[3] , \BUS_ADDR_INTERNAL[2] , \BUS_ADDR_INTERNAL[3] , 
            \BUS_ADDR_INTERNAL[4] , \BUS_ADDR_INTERNAL[5] , \BUS_ADDR_INTERNAL[6] , 
            \BUS_ADDR_INTERNAL[7] , \BUS_ADDR_INTERNAL[13] , \BUS_ADDR_INTERNAL[14] , 
            \BUS_ADDR_INTERNAL[15] , \BUS_ADDR_INTERNAL[16] , \BUS_ADDR_INTERNAL[17] , 
            \BUS_data[4] , \BUS_data[5] , \BUS_data[6] , \BUS_data[7] , 
            \writeData[4] , \writeData[5] , \writeData[6] , \writeData[7] , 
            PIC_DATA_IN_out_2, PIC_DATA_IN_out_1, PIC_DATA_IN_out_4, PIC_DATA_IN_out_3, 
            PIC_DATA_IN_out_6, PIC_DATA_IN_out_5, n18264, lastAddress_31__N_1310, 
            n18271, n18277, n18266, n18262, n18274, n18265, n18276, 
            n17409, n18275, n17423, n18263, n18261, n17275, \BUS_DATA_INTERNAL[1] , 
            \BUS_DATA_INTERNAL[2] , \BUS_DATA_INTERNAL[3] );
    input PIC_DATA_IN_out_7;
    input \BUS_currGrantID[1] ;
    input \BUS_currGrantID[0] ;
    output \BUS_ADDR_INTERNAL[11] ;
    input n18273;
    output \BUS_ADDR_INTERNAL[12] ;
    input n18272;
    input GND_net;
    output [15:0]writeData;
    input LOGIC_CLOCK;
    input PIC_DATA_IN_out_15;
    input PIC_DATA_IN_out_14;
    input PIC_DATA_IN_out_13;
    input PIC_DATA_IN_out_12;
    input PIC_DATA_IN_out_11;
    output \BUS_ADDR_INTERNAL[9] ;
    input n18268;
    output \BUS_ADDR_INTERNAL[10] ;
    input n18269;
    output \BUS_ADDR_INTERNAL[8] ;
    input n18267;
    output OUT_ENABLE;
    input n9950;
    output \PIC_data[0] ;
    output \writeData[10] ;
    input PIC_DATA_IN_out_10;
    output \writeData[9] ;
    input PIC_DATA_IN_out_9;
    output \writeData[8] ;
    input PIC_DATA_IN_out_8;
    input n17298;
    input n17337;
    input n17325;
    input n15534;
    output [7:0]state;
    input n17270;
    input PIC_WE_IN_c;
    input \BUS_data[0] ;
    output \BUS_ADDR_INTERNAL[0] ;
    input PIC_ADDR_IN_c_0;
    output \BUS_ADDR_INTERNAL[1] ;
    input \BUS_ADDR_INTERNAL[1]_adj_1 ;
    output n17384;
    output \BUS_req[2] ;
    output \BUS_ADDR_INTERNAL[18] ;
    input n2642;
    output LOGIC_CLOCK_enable_52;
    input n2504;
    output n17279;
    input PIC_DATA_IN_out_0;
    output WRITE_DONE;
    input n18280;
    input PIC_ADDR_IN_c_1;
    input PIC_ADDR_IN_c_2;
    input PIC_ADDR_IN_c_3;
    input PIC_ADDR_IN_c_4;
    input PIC_ADDR_IN_c_5;
    input PIC_ADDR_IN_c_6;
    input PIC_ADDR_IN_c_7;
    input PIC_ADDR_IN_c_8;
    input PIC_ADDR_IN_c_9;
    input PIC_ADDR_IN_c_10;
    input PIC_ADDR_IN_c_11;
    input PIC_ADDR_IN_c_12;
    input PIC_ADDR_IN_c_13;
    input PIC_ADDR_IN_c_14;
    input PIC_ADDR_IN_c_15;
    input PIC_ADDR_IN_c_16;
    input PIC_ADDR_IN_c_17;
    input PIC_ADDR_IN_c_18;
    input n14;
    output n17434;
    output BUS_DIRECTION_INTERNAL;
    input n18260;
    input n16456;
    input n17276;
    output LOGIC_CLOCK_N_57_enable_3;
    input n17457;
    input n17278;
    output n15571;
    input PIC_OE_c;
    input n15469;
    output PIC_READY_c;
    input [7:0]SpriteRead_yInSprite;
    input \currSprite_size[6] ;
    input \currSprite_size[4] ;
    input \currSprite_size[2] ;
    input n17394;
    output \Sprite_readAddr_13__N_752[0] ;
    output \Sprite_readAddr_13__N_752[2] ;
    output \Sprite_readAddr_13__N_752[3] ;
    output \Sprite_readAddr_13__N_752[4] ;
    output \Sprite_readAddr_13__N_752[6] ;
    output \Sprite_readAddr_13__N_752[5] ;
    output \Sprite_readAddr_13__N_752[8] ;
    output \Sprite_readAddr_13__N_752[7] ;
    output \Sprite_readAddr_13__N_752[10] ;
    output \Sprite_readAddr_13__N_752[9] ;
    output \Sprite_readAddr_13__N_752[12] ;
    output \Sprite_readAddr_13__N_752[11] ;
    output \Sprite_readAddr_13__N_752[13] ;
    input \currSprite_size[1] ;
    output \Sprite_readAddr_13__N_752[1] ;
    input \currSprite_size[3] ;
    input \currSprite_size[5] ;
    input \currSprite_size[7] ;
    input \BUS_data[1] ;
    input \BUS_data[2] ;
    input \BUS_data[3] ;
    output \BUS_ADDR_INTERNAL[2] ;
    output \BUS_ADDR_INTERNAL[3] ;
    output \BUS_ADDR_INTERNAL[4] ;
    output \BUS_ADDR_INTERNAL[5] ;
    output \BUS_ADDR_INTERNAL[6] ;
    output \BUS_ADDR_INTERNAL[7] ;
    output \BUS_ADDR_INTERNAL[13] ;
    output \BUS_ADDR_INTERNAL[14] ;
    output \BUS_ADDR_INTERNAL[15] ;
    output \BUS_ADDR_INTERNAL[16] ;
    output \BUS_ADDR_INTERNAL[17] ;
    input \BUS_data[4] ;
    input \BUS_data[5] ;
    input \BUS_data[6] ;
    input \BUS_data[7] ;
    output \writeData[4] ;
    output \writeData[5] ;
    output \writeData[6] ;
    output \writeData[7] ;
    input PIC_DATA_IN_out_2;
    input PIC_DATA_IN_out_1;
    input PIC_DATA_IN_out_4;
    input PIC_DATA_IN_out_3;
    input PIC_DATA_IN_out_6;
    input PIC_DATA_IN_out_5;
    input n18264;
    input lastAddress_31__N_1310;
    input n18271;
    input n18277;
    input n18266;
    input n18262;
    input n18274;
    input n18265;
    input n18276;
    input n17409;
    input n18275;
    input n17423;
    input n18263;
    input n18261;
    input n17275;
    output \BUS_DATA_INTERNAL[1] ;
    output \BUS_DATA_INTERNAL[2] ;
    output \BUS_DATA_INTERNAL[3] ;
    
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire BUS_DIRECTION_INTERNAL_N_1547 /* synthesis is_clock=1, SET_AS_NETWORK=\PIC_BUS_INTERFACE/BUS_DIRECTION_INTERNAL_N_1547 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(38[8:30])
    wire [16:0]rModDataWrite;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(54[8:21])
    
    wire n15, n5868;
    wire [15:0]writeData_15__N_1719;
    
    wire n14172, n14173, mult_8u_9u_0_cin_lr_0, mult_8u_8u_0_cin_lr_0, 
        LOGIC_CLOCK_enable_248, n7202, n14171;
    wire [15:0]readData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(45[8:16])
    wire [15:0]writeData_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(46[8:17])
    wire [3:0]transferMode;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(50[8:20])
    
    wire n63, n17350, n15491, n8;
    wire [7:0]state_7__N_1600;
    
    wire n15336, n17389, n15335, n15350, LOGIC_CLOCK_enable_216, LOGIC_CLOCK_enable_259;
    wire [7:0]rModDataRead;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(53[8:20])
    
    wire LOGIC_CLOCK_enable_241, BUS_REQ_N_1761, mult_8u_8u_0_cin_lr_0_adj_1773;
    wire [7:0]state_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    wire [7:0]rModDataTrans;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(56[8:21])
    wire [15:0]data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(44[8:12])
    wire [18:0]lastAddress;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(41[8:19])
    
    wire transferMode_3__N_1665, n17390, n17475, n17290, n6, LOGIC_CLOCK_enable_44, 
        n18, n17400, n17364, n15494, n14_adj_1774, n10, BUS_VALID_N_1668, 
        n2780, n16942, n17444, BUS_DIRECTION_INTERNAL_N_1550, n17292, 
        n15460, n9, n17445, n17401, n17352, n17363, LOGIC_CLOCK_enable_249, 
        LOGIC_CLOCK_enable_250, n17474, LOGIC_CLOCK_enable_80;
    wire [9:0]rModDataWrite_15__N_1670;
    
    wire mult_8u_9u_0_pp_3_6, mult_8u_9u_0_pp_2_4, mult_8u_9u_0_pp_1_2;
    wire [16:0]rModDataWrite_15__N_1620;
    
    wire mult_8u_9u_0_cin_lr_2, mult_8u_9u_0_cin_lr_4, mult_8u_9u_0_cin_lr_6, 
        co_mult_8u_9u_0_0_1, mult_8u_9u_0_pp_0_2, co_mult_8u_9u_0_0_2, 
        s_mult_8u_9u_0_0_4, mult_8u_9u_0_pp_0_4, mult_8u_9u_0_pp_0_3, 
        mult_8u_9u_0_pp_1_4, mult_8u_9u_0_pp_1_3, co_mult_8u_9u_0_0_3, 
        s_mult_8u_9u_0_0_5, s_mult_8u_9u_0_0_6, mult_8u_9u_0_pp_0_6, mult_8u_9u_0_pp_0_5, 
        mult_8u_9u_0_pp_1_6, mult_8u_9u_0_pp_1_5, co_mult_8u_9u_0_0_4, 
        s_mult_8u_9u_0_0_7, s_mult_8u_9u_0_0_8, mult_8u_9u_0_pp_0_8, mult_8u_9u_0_pp_0_7, 
        mult_8u_9u_0_pp_1_8, mult_8u_9u_0_pp_1_7, co_mult_8u_9u_0_0_5, 
        s_mult_8u_9u_0_0_9, s_mult_8u_9u_0_0_10, mult_8u_9u_0_pp_0_10, 
        mult_8u_9u_0_pp_0_9, mult_8u_9u_0_pp_1_10, mult_8u_9u_0_pp_1_9, 
        co_mult_8u_9u_0_0_6, s_mult_8u_9u_0_0_11, s_mult_8u_9u_0_0_12, 
        mult_8u_9u_0_pp_1_12, mult_8u_9u_0_pp_1_11, s_mult_8u_9u_0_0_13, 
        co_mult_8u_9u_0_1_1, s_mult_8u_9u_0_1_6, mult_8u_9u_0_pp_2_6, 
        co_mult_8u_9u_0_1_2, s_mult_8u_9u_0_1_7, s_mult_8u_9u_0_1_8, mult_8u_9u_0_pp_2_8, 
        mult_8u_9u_0_pp_2_7, mult_8u_9u_0_pp_3_8, mult_8u_9u_0_pp_3_7, 
        co_mult_8u_9u_0_1_3, s_mult_8u_9u_0_1_9, s_mult_8u_9u_0_1_10, 
        mult_8u_9u_0_pp_2_10, mult_8u_9u_0_pp_2_9, mult_8u_9u_0_pp_3_10, 
        mult_8u_9u_0_pp_3_9, co_mult_8u_9u_0_1_4, s_mult_8u_9u_0_1_11, 
        s_mult_8u_9u_0_1_12, mult_8u_9u_0_pp_2_12, mult_8u_9u_0_pp_2_11, 
        mult_8u_9u_0_pp_3_12, mult_8u_9u_0_pp_3_11, co_mult_8u_9u_0_1_5, 
        s_mult_8u_9u_0_1_13, s_mult_8u_9u_0_1_14, mult_8u_9u_0_pp_2_14, 
        mult_8u_9u_0_pp_2_13, mult_8u_9u_0_pp_3_14, mult_8u_9u_0_pp_3_13, 
        s_mult_8u_9u_0_1_15, s_mult_8u_9u_0_1_16, mult_8u_9u_0_pp_3_16, 
        mult_8u_9u_0_pp_3_15, co_t_mult_8u_9u_0_2_1, co_t_mult_8u_9u_0_2_2, 
        mult_8u_9u_0_pp_2_5, co_t_mult_8u_9u_0_2_3, co_t_mult_8u_9u_0_2_4, 
        co_t_mult_8u_9u_0_2_5, co_t_mult_8u_9u_0_2_6, mco, mco_1, mco_2, 
        mco_3, mco_4, mco_5, mco_6, mco_7, mco_8, mco_9, mco_10, 
        mco_11, mco_12, mco_13, mco_14, mco_15, mult_8u_8u_0_pp_3_6, 
        mult_8u_8u_0_pp_2_4, mult_8u_8u_0_pp_1_2, mult_8u_8u_0_pp_0_9, 
        mfco, mult_8u_8u_0_cin_lr_2, mult_8u_8u_0_pp_1_11, mfco_1, mult_8u_8u_0_cin_lr_4, 
        mult_8u_8u_0_pp_2_13, mfco_2, mult_8u_8u_0_cin_lr_6, co_mult_8u_8u_0_0_1, 
        mult_8u_8u_0_pp_0_2, co_mult_8u_8u_0_0_2, s_mult_8u_8u_0_0_4, 
        mult_8u_8u_0_pp_0_4, mult_8u_8u_0_pp_0_3, mult_8u_8u_0_pp_1_4, 
        mult_8u_8u_0_pp_1_3, co_mult_8u_8u_0_0_3, s_mult_8u_8u_0_0_5, 
        s_mult_8u_8u_0_0_6, mult_8u_8u_0_pp_0_6, mult_8u_8u_0_pp_0_5, 
        mult_8u_8u_0_pp_1_6, mult_8u_8u_0_pp_1_5, co_mult_8u_8u_0_0_4, 
        s_mult_8u_8u_0_0_7, s_mult_8u_8u_0_0_8, mult_8u_8u_0_pp_0_8, mult_8u_8u_0_pp_0_7, 
        mult_8u_8u_0_pp_1_8, mult_8u_8u_0_pp_1_7, co_mult_8u_8u_0_0_5, 
        s_mult_8u_8u_0_0_9, s_mult_8u_8u_0_0_10, mult_8u_8u_0_pp_1_10, 
        mult_8u_8u_0_pp_1_9, co_mult_8u_8u_0_0_6, s_mult_8u_8u_0_0_11, 
        s_mult_8u_8u_0_0_12, s_mult_8u_8u_0_0_13, co_mult_8u_8u_0_1_1, 
        s_mult_8u_8u_0_1_6, mult_8u_8u_0_pp_2_6, co_mult_8u_8u_0_1_2, 
        s_mult_8u_8u_0_1_7, s_mult_8u_8u_0_1_8, mult_8u_8u_0_pp_2_8, mult_8u_8u_0_pp_2_7, 
        mult_8u_8u_0_pp_3_8, mult_8u_8u_0_pp_3_7, co_mult_8u_8u_0_1_3, 
        s_mult_8u_8u_0_1_9, s_mult_8u_8u_0_1_10, mult_8u_8u_0_pp_2_10, 
        mult_8u_8u_0_pp_2_9, mult_8u_8u_0_pp_3_10, mult_8u_8u_0_pp_3_9, 
        co_mult_8u_8u_0_1_4, s_mult_8u_8u_0_1_11, s_mult_8u_8u_0_1_12, 
        mult_8u_8u_0_pp_2_12, mult_8u_8u_0_pp_2_11, mult_8u_8u_0_pp_3_12, 
        mult_8u_8u_0_pp_3_11, s_mult_8u_8u_0_1_13, s_mult_8u_8u_0_1_14, 
        mult_8u_8u_0_pp_3_14, mult_8u_8u_0_pp_3_13, co_t_mult_8u_8u_0_2_1, 
        co_t_mult_8u_8u_0_2_2, mult_8u_8u_0_pp_2_5, co_t_mult_8u_8u_0_2_3, 
        co_t_mult_8u_8u_0_2_4, co_t_mult_8u_8u_0_2_5, mco_adj_1775, mco_1_adj_1776, 
        mco_2_adj_1777, mco_3_adj_1778, mco_4_adj_1779, mco_5_adj_1780, 
        mco_6_adj_1781, mco_7_adj_1782, mco_8_adj_1783, mco_9_adj_1784, 
        mco_10_adj_1785, mco_11_adj_1786, n14117, n14116, n14115, 
        n14114, mult_8u_8u_0_pp_3_6_adj_1787, mult_8u_8u_0_pp_2_4_adj_1788, 
        mult_8u_8u_0_pp_1_2_adj_1789;
    wire [15:0]rModDataWrite_15__N_1637;
    
    wire mult_8u_8u_0_pp_0_9_adj_1790, mfco_adj_1791, mult_8u_8u_0_cin_lr_2_adj_1792, 
        mult_8u_8u_0_pp_1_11_adj_1793, mfco_1_adj_1794, mult_8u_8u_0_cin_lr_4_adj_1795, 
        mult_8u_8u_0_pp_2_13_adj_1796, mfco_2_adj_1797, mult_8u_8u_0_cin_lr_6_adj_1798, 
        mult_8u_8u_0_pp_3_15, mfco_3, co_mult_8u_8u_0_0_1_adj_1799, mult_8u_8u_0_pp_0_2_adj_1800, 
        co_mult_8u_8u_0_0_2_adj_1801, s_mult_8u_8u_0_0_4_adj_1802, mult_8u_8u_0_pp_0_4_adj_1803, 
        mult_8u_8u_0_pp_0_3_adj_1804, mult_8u_8u_0_pp_1_4_adj_1805, mult_8u_8u_0_pp_1_3_adj_1806, 
        co_mult_8u_8u_0_0_3_adj_1807, s_mult_8u_8u_0_0_5_adj_1808, s_mult_8u_8u_0_0_6_adj_1809, 
        mult_8u_8u_0_pp_0_6_adj_1810, mult_8u_8u_0_pp_0_5_adj_1811, mult_8u_8u_0_pp_1_6_adj_1812, 
        mult_8u_8u_0_pp_1_5_adj_1813, co_mult_8u_8u_0_0_4_adj_1814, s_mult_8u_8u_0_0_7_adj_1815, 
        s_mult_8u_8u_0_0_8_adj_1816, mult_8u_8u_0_pp_0_8_adj_1817, mult_8u_8u_0_pp_0_7_adj_1818, 
        mult_8u_8u_0_pp_1_8_adj_1819, mult_8u_8u_0_pp_1_7_adj_1820, co_mult_8u_8u_0_0_5_adj_1821, 
        s_mult_8u_8u_0_0_9_adj_1822, s_mult_8u_8u_0_0_10_adj_1823, mult_8u_8u_0_pp_1_10_adj_1824, 
        mult_8u_8u_0_pp_1_9_adj_1825, co_mult_8u_8u_0_0_6_adj_1826, s_mult_8u_8u_0_0_11_adj_1827, 
        s_mult_8u_8u_0_0_12_adj_1828, s_mult_8u_8u_0_0_13_adj_1829, co_mult_8u_8u_0_1_1_adj_1830, 
        s_mult_8u_8u_0_1_6_adj_1831, mult_8u_8u_0_pp_2_6_adj_1832, co_mult_8u_8u_0_1_2_adj_1833, 
        s_mult_8u_8u_0_1_7_adj_1834, s_mult_8u_8u_0_1_8_adj_1835, mult_8u_8u_0_pp_2_8_adj_1836, 
        mult_8u_8u_0_pp_2_7_adj_1837, mult_8u_8u_0_pp_3_8_adj_1838, mult_8u_8u_0_pp_3_7_adj_1839, 
        co_mult_8u_8u_0_1_3_adj_1840, s_mult_8u_8u_0_1_9_adj_1841, s_mult_8u_8u_0_1_10_adj_1842, 
        mult_8u_8u_0_pp_2_10_adj_1843, mult_8u_8u_0_pp_2_9_adj_1844, mult_8u_8u_0_pp_3_10_adj_1845, 
        mult_8u_8u_0_pp_3_9_adj_1846, co_mult_8u_8u_0_1_4_adj_1847, s_mult_8u_8u_0_1_11_adj_1848, 
        s_mult_8u_8u_0_1_12_adj_1849, mult_8u_8u_0_pp_2_12_adj_1850, mult_8u_8u_0_pp_2_11_adj_1851, 
        mult_8u_8u_0_pp_3_12_adj_1852, mult_8u_8u_0_pp_3_11_adj_1853, co_mult_8u_8u_0_1_5, 
        s_mult_8u_8u_0_1_13_adj_1854, s_mult_8u_8u_0_1_14_adj_1855, mult_8u_8u_0_pp_3_14_adj_1856, 
        mult_8u_8u_0_pp_3_13_adj_1857, s_mult_8u_8u_0_1_15, co_t_mult_8u_8u_0_2_1_adj_1858, 
        co_t_mult_8u_8u_0_2_2_adj_1859, mult_8u_8u_0_pp_2_5_adj_1860, co_t_mult_8u_8u_0_2_3_adj_1861, 
        co_t_mult_8u_8u_0_2_4_adj_1862, co_t_mult_8u_8u_0_2_5_adj_1863, 
        co_t_mult_8u_8u_0_2_6, mco_adj_1864, mco_1_adj_1865, mco_2_adj_1866, 
        mco_3_adj_1867, mco_4_adj_1868, mco_5_adj_1869, mco_6_adj_1870, 
        mco_7_adj_1871, mco_8_adj_1872, mco_9_adj_1873, mco_10_adj_1874, 
        mco_11_adj_1875, n9_adj_1876, n14_adj_1877, n10_adj_1878, LOGIC_CLOCK_enable_251, 
        LOGIC_CLOCK_enable_252, n14103, n14102, n14101, n14100, n14099, 
        n14098, n14097, n14289, n14288, n14287, n14286, n14285, 
        n14284, n14283, n14282, n14281, n14280, n14279, n6105, 
        n15454, n13663, n13667, n13666, n15599, n16943, n13665, 
        n15657, n17324, n15495, n15490, n14177, n14176, n14175, 
        n14174, n16941, n13664, n15577, n12, n6_adj_1879;
    
    LUT4 mux_725_i8_4_lut (.A(rModDataWrite[15]), .B(PIC_DATA_IN_out_7), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i8_4_lut.init = 16'h0aca;
    CCU2D add_10511_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n18273), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n18272), 
          .CIN(n14172), .COUT(n14173));
    defparam add_10511_5.INIT0 = 16'h00ce;
    defparam add_10511_5.INIT1 = 16'h00ce;
    defparam add_10511_5.INJECT1_0 = "NO";
    defparam add_10511_5.INJECT1_1 = "NO";
    FADD2B mult_8u_9u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_8u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FD1P3IX writeData_i0_i15 (.D(PIC_DATA_IN_out_15), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(writeData[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i15.GSR = "DISABLED";
    FD1P3IX writeData_i0_i14 (.D(PIC_DATA_IN_out_14), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(writeData[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i14.GSR = "DISABLED";
    FD1P3IX writeData_i0_i13 (.D(PIC_DATA_IN_out_13), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(writeData[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i13.GSR = "DISABLED";
    FD1P3IX writeData_i0_i12 (.D(PIC_DATA_IN_out_12), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(writeData[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i12.GSR = "DISABLED";
    FD1P3IX writeData_i0_i11 (.D(PIC_DATA_IN_out_11), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(writeData[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i11.GSR = "DISABLED";
    CCU2D add_10511_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[9] ), .D0(n18268), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n18269), 
          .CIN(n14171), .COUT(n14172));
    defparam add_10511_3.INIT0 = 16'h00ce;
    defparam add_10511_3.INIT1 = 16'hff31;
    defparam add_10511_3.INJECT1_0 = "NO";
    defparam add_10511_3.INJECT1_1 = "NO";
    CCU2D add_10511_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), 
          .D1(n18267), .COUT(n14171));
    defparam add_10511_1.INIT0 = 16'hF000;
    defparam add_10511_1.INIT1 = 16'h00ce;
    defparam add_10511_1.INJECT1_0 = "NO";
    defparam add_10511_1.INJECT1_1 = "NO";
    LUT4 i6615_4_lut (.A(readData[0]), .B(OUT_ENABLE), .C(writeData_c[0]), 
         .D(n9950), .Z(\PIC_data[0] )) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(66[18:70])
    defparam i6615_4_lut.init = 16'h88c0;
    FD1P3IX writeData_i0_i10 (.D(PIC_DATA_IN_out_10), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(\writeData[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i10.GSR = "DISABLED";
    FD1P3IX writeData_i0_i9 (.D(PIC_DATA_IN_out_9), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(\writeData[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i9.GSR = "DISABLED";
    FD1P3IX writeData_i0_i8 (.D(PIC_DATA_IN_out_8), .SP(LOGIC_CLOCK_enable_248), 
            .CD(n7202), .CK(LOGIC_CLOCK), .Q(\writeData[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i8.GSR = "DISABLED";
    LUT4 i6606_2_lut (.A(transferMode[0]), .B(n63), .Z(readData[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(76[2] 77[32])
    defparam i6606_2_lut.init = 16'h2222;
    LUT4 i3_4_lut (.A(n17298), .B(n17337), .C(n17325), .D(n15534), .Z(n63)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(76[58:69])
    defparam i3_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut (.A(state[1]), .B(n17350), .C(n15491), .D(n8), .Z(state_7__N_1600[1])) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcec;
    LUT4 i2_4_lut (.A(n15336), .B(n17389), .C(n17270), .D(state[4]), 
         .Z(n8)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    defparam i2_4_lut.init = 16'h3022;
    LUT4 i2_3_lut (.A(n15335), .B(PIC_WE_IN_c), .C(n15350), .Z(n15336)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    FD1P3AX transferMode_i0_i0 (.D(\BUS_data[0] ), .SP(LOGIC_CLOCK_enable_216), 
            .CK(LOGIC_CLOCK), .Q(transferMode[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i0.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i1 (.D(PIC_ADDR_IN_c_0), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i1.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i0 (.D(\BUS_data[0] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i0.GSR = "DISABLED";
    LUT4 PIC_addr_31__I_0_i2_2_lut_rep_376_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[1] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(\BUS_ADDR_INTERNAL[1]_adj_1 ), 
         .Z(n17384)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam PIC_addr_31__I_0_i2_2_lut_rep_376_3_lut_4_lut_4_lut.init = 16'h2c20;
    FD1S3DX BUS_REQ_266 (.D(BUS_REQ_N_1761), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_1547), 
            .Q(\BUS_req[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_REQ_266.GSR = "DISABLED";
    FADD2B mult_8u_8u_0_cin_lr_add_0_adj_210 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_0_adj_1773)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FD1P3AX writeData_i0_i0 (.D(writeData_15__N_1719[0]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(writeData_c[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i0.GSR = "DISABLED";
    FD1S3DX state_i0 (.D(state_7__N_1600[0]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_1547), 
            .Q(state_c[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i0.GSR = "DISABLED";
    LUT4 BUS_VALID_N_450_I_0_2_lut_rep_280_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[18] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(n2642), 
         .Z(LOGIC_CLOCK_enable_52)) /* synthesis lut_function=(!(A (B+(D))+!A (B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam BUS_VALID_N_450_I_0_2_lut_rep_280_3_lut_4_lut_4_lut.init = 16'h0023;
    FD1P3AX rModDataTrans_i0_i0 (.D(data[8]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i0.GSR = "DISABLED";
    LUT4 i13105_2_lut_rep_271_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[18] ), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(n2504), 
         .Z(n17279)) /* synthesis lut_function=(A (B+(D))+!A (B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i13105_2_lut_rep_271_3_lut_4_lut_4_lut.init = 16'hffdc;
    FD1S1A PIC_ADDR_IN_18__I_0_i1 (.D(PIC_ADDR_IN_c_0), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i1.GSR = "DISABLED";
    LUT4 mux_725_i1_4_lut (.A(rModDataWrite[8]), .B(PIC_DATA_IN_out_0), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i1_4_lut.init = 16'h0aca;
    FD1S3DX WRITE_DONE_264 (.D(n18280), .CK(LOGIC_CLOCK), .CD(transferMode_3__N_1665), 
            .Q(WRITE_DONE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam WRITE_DONE_264.GSR = "DISABLED";
    LUT4 i6874_2_lut (.A(PIC_DATA_IN_out_8), .B(PIC_WE_IN_c), .Z(data[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6874_2_lut.init = 16'h2222;
    FD1S1A PIC_ADDR_IN_18__I_0_i2 (.D(PIC_ADDR_IN_c_1), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i2.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i3 (.D(PIC_ADDR_IN_c_2), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i3.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i4 (.D(PIC_ADDR_IN_c_3), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i4.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i5 (.D(PIC_ADDR_IN_c_4), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i5.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i6 (.D(PIC_ADDR_IN_c_5), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i6.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i7 (.D(PIC_ADDR_IN_c_6), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i7.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i8 (.D(PIC_ADDR_IN_c_7), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i8.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i9 (.D(PIC_ADDR_IN_c_8), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i9.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i10 (.D(PIC_ADDR_IN_c_9), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i10.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i11 (.D(PIC_ADDR_IN_c_10), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i11.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i12 (.D(PIC_ADDR_IN_c_11), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i12.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i13 (.D(PIC_ADDR_IN_c_12), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i13.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i14 (.D(PIC_ADDR_IN_c_13), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i14.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i15 (.D(PIC_ADDR_IN_c_14), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i15.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i16 (.D(PIC_ADDR_IN_c_15), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i16.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i17 (.D(PIC_ADDR_IN_c_16), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[16])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i17.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i18 (.D(PIC_ADDR_IN_c_17), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[17])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i18.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i19 (.D(PIC_ADDR_IN_c_18), .CK(BUS_DIRECTION_INTERNAL_N_1547), 
           .Q(lastAddress[18])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i19.GSR = "DISABLED";
    LUT4 i7955_3_lut_4_lut_then_4_lut (.A(n17390), .B(n14), .C(state_c[2]), 
         .D(state[1]), .Z(n17475)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    defparam i7955_3_lut_4_lut_then_4_lut.init = 16'hfffb;
    LUT4 i4_4_lut (.A(n17290), .B(n14), .C(state[1]), .D(n6), .Z(LOGIC_CLOCK_enable_44)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0800;
    LUT4 i13039_4_lut (.A(state_c[0]), .B(n18), .C(n17400), .D(n17364), 
         .Z(n15494)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i13039_4_lut.init = 16'h0002;
    LUT4 i1_3_lut (.A(PIC_WE_IN_c), .B(n15350), .C(n15335), .Z(n18)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i1_3_lut.init = 16'h5454;
    LUT4 i7_4_lut (.A(PIC_DATA_IN_out_8), .B(n14_adj_1774), .C(n10), .D(PIC_DATA_IN_out_14), 
         .Z(n15350)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(PIC_DATA_IN_out_11), .B(PIC_DATA_IN_out_9), .C(PIC_DATA_IN_out_13), 
         .D(PIC_DATA_IN_out_15), .Z(n14_adj_1774)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i2_2_lut (.A(PIC_DATA_IN_out_10), .B(PIC_DATA_IN_out_12), .Z(n10)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_211 (.A(transferMode[2]), .B(transferMode[3]), .C(transferMode[1]), 
         .D(transferMode[0]), .Z(n15335)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_211.init = 16'hfeff;
    LUT4 i2_2_lut_rep_426 (.A(state_c[2]), .B(state_c[0]), .Z(n17434)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i2_2_lut_rep_426.init = 16'h4444;
    FD1P3AX BUS_DIRECTION_INTERNAL_272 (.D(n15494), .SP(LOGIC_CLOCK_enable_44), 
            .CK(LOGIC_CLOCK), .Q(BUS_DIRECTION_INTERNAL)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_DIRECTION_INTERNAL_272.GSR = "DISABLED";
    LUT4 transferMode_3__I_197_2_lut_3_lut (.A(BUS_VALID_N_1668), .B(n2780), 
         .C(n18260), .Z(transferMode_3__N_1665)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam transferMode_3__I_197_2_lut_3_lut.init = 16'hfdfd;
    LUT4 i13074_3_lut_4_lut (.A(BUS_VALID_N_1668), .B(n2780), .C(n16456), 
         .D(n17276), .Z(LOGIC_CLOCK_N_57_enable_3)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam i13074_3_lut_4_lut.init = 16'hd000;
    LUT4 OUT_ENABLE_I_0_3_lut_4_lut (.A(BUS_VALID_N_1668), .B(n2780), .C(n18260), 
         .D(n17457), .Z(OUT_ENABLE)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam OUT_ENABLE_I_0_3_lut_4_lut.init = 16'h202f;
    LUT4 i11917_3_lut_4_lut (.A(BUS_VALID_N_1668), .B(n2780), .C(n17278), 
         .D(n18260), .Z(n15571)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam i11917_3_lut_4_lut.init = 16'hf200;
    LUT4 n6241_bdd_2_lut_13374_4_lut (.A(n17434), .B(n15336), .C(n17390), 
         .D(state[4]), .Z(n16942)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam n6241_bdd_2_lut_13374_4_lut.init = 16'hff02;
    LUT4 i2_3_lut_4_lut (.A(n17364), .B(n17400), .C(PIC_WE_IN_c), .D(state_c[0]), 
         .Z(n5868)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_282_3_lut_4_lut (.A(PIC_OE_c), .B(PIC_WE_IN_c), .C(n17444), 
         .D(BUS_DIRECTION_INTERNAL_N_1550), .Z(n17290)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam i1_2_lut_rep_282_3_lut_4_lut.init = 16'h0700;
    LUT4 i1_2_lut_rep_284_3_lut (.A(PIC_OE_c), .B(PIC_WE_IN_c), .C(BUS_DIRECTION_INTERNAL_N_1550), 
         .Z(n17292)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam i1_2_lut_rep_284_3_lut.init = 16'h7070;
    LUT4 BUS_DIRECTION_INTERNAL_I_194_2_lut_3_lut (.A(PIC_OE_c), .B(PIC_WE_IN_c), 
         .C(BUS_DIRECTION_INTERNAL_N_1550), .Z(BUS_DIRECTION_INTERNAL_N_1547)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam BUS_DIRECTION_INTERNAL_I_194_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i3_2_lut_3_lut_4_lut (.A(PIC_OE_c), .B(PIC_WE_IN_c), .C(n15460), 
         .D(BUS_DIRECTION_INTERNAL_N_1550), .Z(n9)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam i3_2_lut_3_lut_4_lut.init = 16'h7000;
    LUT4 i1_2_lut_rep_436 (.A(state_c[2]), .B(state_c[3]), .Z(n17444)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_436.init = 16'heeee;
    LUT4 i1_2_lut_rep_392_3_lut (.A(state_c[2]), .B(state_c[3]), .C(state[1]), 
         .Z(n17400)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_392_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_381_3_lut_4_lut (.A(state_c[2]), .B(state_c[3]), .C(n17445), 
         .D(state_c[5]), .Z(n17389)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_381_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_437 (.A(state_c[6]), .B(state_c[7]), .Z(n17445)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_437.init = 16'heeee;
    LUT4 i2_3_lut_rep_382_4_lut (.A(state_c[6]), .B(state_c[7]), .C(state_c[3]), 
         .D(state_c[5]), .Z(n17390)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_382_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_393_3_lut (.A(state_c[6]), .B(state_c[7]), .C(state_c[5]), 
         .Z(n17401)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_393_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(state_c[6]), .B(state_c[7]), .C(state[4]), 
         .D(state_c[5]), .Z(n17352)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_355_3_lut_4_lut (.A(state_c[6]), .B(state_c[7]), .C(state[4]), 
         .D(state_c[5]), .Z(n17363)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_355_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_356_3_lut_4_lut (.A(state_c[6]), .B(state_c[7]), .C(state[4]), 
         .D(state_c[5]), .Z(n17364)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_356_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_212 (.A(n15460), .B(n17350), .C(n17270), .D(state_c[2]), 
         .Z(LOGIC_CLOCK_enable_249)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_212.init = 16'hcecc;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state_c[6]), .B(state_c[7]), .C(state_c[0]), 
         .D(state_c[5]), .Z(n6)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_213 (.A(n15469), .B(n17350), .C(n17352), .D(state_c[3]), 
         .Z(LOGIC_CLOCK_enable_250)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_213.init = 16'heccc;
    LUT4 i7955_3_lut_4_lut_else_4_lut (.A(n17401), .B(state_c[2]), .C(state_c[3]), 
         .Z(n17474)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    defparam i7955_3_lut_4_lut_else_4_lut.init = 16'h0101;
    FD1P3DX PIC_READY_267 (.D(n18280), .SP(LOGIC_CLOCK_enable_80), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_1547), .Q(PIC_READY_c)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam PIC_READY_267.GSR = "DISABLED";
    AND2 AND2_t0 (.A(rModDataWrite_15__N_1670[0]), .B(rModDataRead[6]), 
         .Z(mult_8u_9u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(134[10:63])
    AND2 AND2_t1 (.A(rModDataWrite_15__N_1670[0]), .B(rModDataRead[4]), 
         .Z(mult_8u_9u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(132[10:63])
    AND2 AND2_t2 (.A(rModDataWrite_15__N_1670[0]), .B(rModDataRead[2]), 
         .Z(mult_8u_9u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(130[10:63])
    AND2 AND2_t3 (.A(rModDataWrite_15__N_1670[0]), .B(rModDataRead[0]), 
         .Z(rModDataWrite_15__N_1620[0])) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(128[10:63])
    FADD2B mult_8u_9u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_mult_8u_9u_0_0_1 (.A0(GND_net), .A1(mult_8u_9u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_8u_9u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_8u_9u_0_0_1), 
           .S1(rModDataWrite_15__N_1620[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_2 (.A0(mult_8u_9u_0_pp_0_3), .A1(mult_8u_9u_0_pp_0_4), 
           .B0(mult_8u_9u_0_pp_1_3), .B1(mult_8u_9u_0_pp_1_4), .CI(co_mult_8u_9u_0_0_1), 
           .COUT(co_mult_8u_9u_0_0_2), .S0(rModDataWrite_15__N_1620[3]), 
           .S1(s_mult_8u_9u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_3 (.A0(mult_8u_9u_0_pp_0_5), .A1(mult_8u_9u_0_pp_0_6), 
           .B0(mult_8u_9u_0_pp_1_5), .B1(mult_8u_9u_0_pp_1_6), .CI(co_mult_8u_9u_0_0_2), 
           .COUT(co_mult_8u_9u_0_0_3), .S0(s_mult_8u_9u_0_0_5), .S1(s_mult_8u_9u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_4 (.A0(mult_8u_9u_0_pp_0_7), .A1(mult_8u_9u_0_pp_0_8), 
           .B0(mult_8u_9u_0_pp_1_7), .B1(mult_8u_9u_0_pp_1_8), .CI(co_mult_8u_9u_0_0_3), 
           .COUT(co_mult_8u_9u_0_0_4), .S0(s_mult_8u_9u_0_0_7), .S1(s_mult_8u_9u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_5 (.A0(mult_8u_9u_0_pp_0_9), .A1(mult_8u_9u_0_pp_0_10), 
           .B0(mult_8u_9u_0_pp_1_9), .B1(mult_8u_9u_0_pp_1_10), .CI(co_mult_8u_9u_0_0_4), 
           .COUT(co_mult_8u_9u_0_0_5), .S0(s_mult_8u_9u_0_0_9), .S1(s_mult_8u_9u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_9u_0_pp_1_11), 
           .B1(mult_8u_9u_0_pp_1_12), .CI(co_mult_8u_9u_0_0_5), .COUT(co_mult_8u_9u_0_0_6), 
           .S0(s_mult_8u_9u_0_0_11), .S1(s_mult_8u_9u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_mult_8u_9u_0_0_7 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_8u_9u_0_0_6), .S0(s_mult_8u_9u_0_0_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_mult_8u_9u_0_1_1 (.A0(GND_net), .A1(mult_8u_9u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_8u_9u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_8u_9u_0_1_1), 
           .S1(s_mult_8u_9u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_2 (.A0(mult_8u_9u_0_pp_2_7), .A1(mult_8u_9u_0_pp_2_8), 
           .B0(mult_8u_9u_0_pp_3_7), .B1(mult_8u_9u_0_pp_3_8), .CI(co_mult_8u_9u_0_1_1), 
           .COUT(co_mult_8u_9u_0_1_2), .S0(s_mult_8u_9u_0_1_7), .S1(s_mult_8u_9u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_3 (.A0(mult_8u_9u_0_pp_2_9), .A1(mult_8u_9u_0_pp_2_10), 
           .B0(mult_8u_9u_0_pp_3_9), .B1(mult_8u_9u_0_pp_3_10), .CI(co_mult_8u_9u_0_1_2), 
           .COUT(co_mult_8u_9u_0_1_3), .S0(s_mult_8u_9u_0_1_9), .S1(s_mult_8u_9u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_4 (.A0(mult_8u_9u_0_pp_2_11), .A1(mult_8u_9u_0_pp_2_12), 
           .B0(mult_8u_9u_0_pp_3_11), .B1(mult_8u_9u_0_pp_3_12), .CI(co_mult_8u_9u_0_1_3), 
           .COUT(co_mult_8u_9u_0_1_4), .S0(s_mult_8u_9u_0_1_11), .S1(s_mult_8u_9u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_5 (.A0(mult_8u_9u_0_pp_2_13), .A1(mult_8u_9u_0_pp_2_14), 
           .B0(mult_8u_9u_0_pp_3_13), .B1(mult_8u_9u_0_pp_3_14), .CI(co_mult_8u_9u_0_1_4), 
           .COUT(co_mult_8u_9u_0_1_5), .S0(s_mult_8u_9u_0_1_13), .S1(s_mult_8u_9u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_9u_0_pp_3_15), 
           .B1(mult_8u_9u_0_pp_3_16), .CI(co_mult_8u_9u_0_1_5), .S0(s_mult_8u_9u_0_1_15), 
           .S1(s_mult_8u_9u_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_t_mult_8u_9u_0_2_1 (.A0(GND_net), .A1(s_mult_8u_9u_0_0_4), 
           .B0(GND_net), .B1(mult_8u_9u_0_pp_2_4), .CI(GND_net), .COUT(co_t_mult_8u_9u_0_2_1), 
           .S1(rModDataWrite_15__N_1620[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_2 (.A0(s_mult_8u_9u_0_0_5), .A1(s_mult_8u_9u_0_0_6), 
           .B0(mult_8u_9u_0_pp_2_5), .B1(s_mult_8u_9u_0_1_6), .CI(co_t_mult_8u_9u_0_2_1), 
           .COUT(co_t_mult_8u_9u_0_2_2), .S0(rModDataWrite_15__N_1620[5]), 
           .S1(rModDataWrite_15__N_1620[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_3 (.A0(s_mult_8u_9u_0_0_7), .A1(s_mult_8u_9u_0_0_8), 
           .B0(s_mult_8u_9u_0_1_7), .B1(s_mult_8u_9u_0_1_8), .CI(co_t_mult_8u_9u_0_2_2), 
           .COUT(co_t_mult_8u_9u_0_2_3), .S0(rModDataWrite_15__N_1620[7]), 
           .S1(rModDataWrite_15__N_1620[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_4 (.A0(s_mult_8u_9u_0_0_9), .A1(s_mult_8u_9u_0_0_10), 
           .B0(s_mult_8u_9u_0_1_9), .B1(s_mult_8u_9u_0_1_10), .CI(co_t_mult_8u_9u_0_2_3), 
           .COUT(co_t_mult_8u_9u_0_2_4), .S0(rModDataWrite_15__N_1620[9]), 
           .S1(rModDataWrite_15__N_1620[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_5 (.A0(s_mult_8u_9u_0_0_11), .A1(s_mult_8u_9u_0_0_12), 
           .B0(s_mult_8u_9u_0_1_11), .B1(s_mult_8u_9u_0_1_12), .CI(co_t_mult_8u_9u_0_2_4), 
           .COUT(co_t_mult_8u_9u_0_2_5), .S0(rModDataWrite_15__N_1620[11]), 
           .S1(rModDataWrite_15__N_1620[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_6 (.A0(s_mult_8u_9u_0_0_13), .A1(GND_net), 
           .B0(s_mult_8u_9u_0_1_13), .B1(s_mult_8u_9u_0_1_14), .CI(co_t_mult_8u_9u_0_2_5), 
           .COUT(co_t_mult_8u_9u_0_2_6), .S0(rModDataWrite_15__N_1620[13]), 
           .S1(rModDataWrite_15__N_1620[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_7 (.A0(GND_net), .A1(GND_net), .B0(s_mult_8u_9u_0_1_15), 
           .B1(s_mult_8u_9u_0_1_16), .CI(co_t_mult_8u_9u_0_2_6), .S0(rModDataWrite_15__N_1620[15])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_0 (.A0(rModDataWrite_15__N_1670[0]), .A1(rModDataWrite_15__N_1670[1]), 
          .A2(rModDataWrite_15__N_1670[1]), .A3(rModDataWrite_15__N_1670[2]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mult_8u_9u_0_cin_lr_0), .CO(mco), 
          .P0(rModDataWrite_15__N_1620[1]), .P1(mult_8u_9u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_1 (.A0(rModDataWrite_15__N_1670[2]), .A1(rModDataWrite_15__N_1670[3]), 
          .A2(rModDataWrite_15__N_1670[3]), .A3(rModDataWrite_15__N_1670[4]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mco), .CO(mco_1), .P0(mult_8u_9u_0_pp_0_3), 
          .P1(mult_8u_9u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_2 (.A0(rModDataWrite_15__N_1670[4]), .A1(rModDataWrite_15__N_1670[5]), 
          .A2(rModDataWrite_15__N_1670[5]), .A3(rModDataWrite_15__N_1670[6]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mco_1), .CO(mco_2), .P0(mult_8u_9u_0_pp_0_5), 
          .P1(mult_8u_9u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_3 (.A0(rModDataWrite_15__N_1670[6]), .A1(rModDataWrite_15__N_1670[7]), 
          .A2(rModDataWrite_15__N_1670[7]), .A3(rModDataWrite_15__N_1670[8]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mco_2), .CO(mco_3), .P0(mult_8u_9u_0_pp_0_7), 
          .P1(mult_8u_9u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_4 (.A0(rModDataWrite_15__N_1670[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[1]), .B1(rModDataRead[0]), 
          .B2(rModDataRead[1]), .B3(rModDataRead[0]), .CI(mco_3), .P0(mult_8u_9u_0_pp_0_9), 
          .P1(mult_8u_9u_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_0 (.A0(rModDataWrite_15__N_1670[0]), .A1(rModDataWrite_15__N_1670[1]), 
          .A2(rModDataWrite_15__N_1670[1]), .A3(rModDataWrite_15__N_1670[2]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mult_8u_9u_0_cin_lr_2), .CO(mco_4), 
          .P0(mult_8u_9u_0_pp_1_3), .P1(mult_8u_9u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_1 (.A0(rModDataWrite_15__N_1670[2]), .A1(rModDataWrite_15__N_1670[3]), 
          .A2(rModDataWrite_15__N_1670[3]), .A3(rModDataWrite_15__N_1670[4]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mco_4), .CO(mco_5), .P0(mult_8u_9u_0_pp_1_5), 
          .P1(mult_8u_9u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_2 (.A0(rModDataWrite_15__N_1670[4]), .A1(rModDataWrite_15__N_1670[5]), 
          .A2(rModDataWrite_15__N_1670[5]), .A3(rModDataWrite_15__N_1670[6]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mco_5), .CO(mco_6), .P0(mult_8u_9u_0_pp_1_7), 
          .P1(mult_8u_9u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_3 (.A0(rModDataWrite_15__N_1670[6]), .A1(rModDataWrite_15__N_1670[7]), 
          .A2(rModDataWrite_15__N_1670[7]), .A3(rModDataWrite_15__N_1670[8]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mco_6), .CO(mco_7), .P0(mult_8u_9u_0_pp_1_9), 
          .P1(mult_8u_9u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_4 (.A0(rModDataWrite_15__N_1670[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[3]), .B1(rModDataRead[2]), 
          .B2(rModDataRead[3]), .B3(rModDataRead[2]), .CI(mco_7), .P0(mult_8u_9u_0_pp_1_11), 
          .P1(mult_8u_9u_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_0 (.A0(rModDataWrite_15__N_1670[0]), .A1(rModDataWrite_15__N_1670[1]), 
          .A2(rModDataWrite_15__N_1670[1]), .A3(rModDataWrite_15__N_1670[2]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mult_8u_9u_0_cin_lr_4), .CO(mco_8), 
          .P0(mult_8u_9u_0_pp_2_5), .P1(mult_8u_9u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_1 (.A0(rModDataWrite_15__N_1670[2]), .A1(rModDataWrite_15__N_1670[3]), 
          .A2(rModDataWrite_15__N_1670[3]), .A3(rModDataWrite_15__N_1670[4]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mco_8), .CO(mco_9), .P0(mult_8u_9u_0_pp_2_7), 
          .P1(mult_8u_9u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_2 (.A0(rModDataWrite_15__N_1670[4]), .A1(rModDataWrite_15__N_1670[5]), 
          .A2(rModDataWrite_15__N_1670[5]), .A3(rModDataWrite_15__N_1670[6]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mco_9), .CO(mco_10), .P0(mult_8u_9u_0_pp_2_9), 
          .P1(mult_8u_9u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_3 (.A0(rModDataWrite_15__N_1670[6]), .A1(rModDataWrite_15__N_1670[7]), 
          .A2(rModDataWrite_15__N_1670[7]), .A3(rModDataWrite_15__N_1670[8]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mco_10), .CO(mco_11), .P0(mult_8u_9u_0_pp_2_11), 
          .P1(mult_8u_9u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_4 (.A0(rModDataWrite_15__N_1670[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[5]), .B1(rModDataRead[4]), 
          .B2(rModDataRead[5]), .B3(rModDataRead[4]), .CI(mco_11), .P0(mult_8u_9u_0_pp_2_13), 
          .P1(mult_8u_9u_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_0 (.A0(rModDataWrite_15__N_1670[0]), .A1(rModDataWrite_15__N_1670[1]), 
          .A2(rModDataWrite_15__N_1670[1]), .A3(rModDataWrite_15__N_1670[2]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mult_8u_9u_0_cin_lr_6), .CO(mco_12), 
          .P0(mult_8u_9u_0_pp_3_7), .P1(mult_8u_9u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_1 (.A0(rModDataWrite_15__N_1670[2]), .A1(rModDataWrite_15__N_1670[3]), 
          .A2(rModDataWrite_15__N_1670[3]), .A3(rModDataWrite_15__N_1670[4]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mco_12), .CO(mco_13), .P0(mult_8u_9u_0_pp_3_9), 
          .P1(mult_8u_9u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_2 (.A0(rModDataWrite_15__N_1670[4]), .A1(rModDataWrite_15__N_1670[5]), 
          .A2(rModDataWrite_15__N_1670[5]), .A3(rModDataWrite_15__N_1670[6]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mco_13), .CO(mco_14), .P0(mult_8u_9u_0_pp_3_11), 
          .P1(mult_8u_9u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_3 (.A0(rModDataWrite_15__N_1670[6]), .A1(rModDataWrite_15__N_1670[7]), 
          .A2(rModDataWrite_15__N_1670[7]), .A3(rModDataWrite_15__N_1670[8]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mco_14), .CO(mco_15), .P0(mult_8u_9u_0_pp_3_13), 
          .P1(mult_8u_9u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_4 (.A0(rModDataWrite_15__N_1670[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[7]), .B1(rModDataRead[6]), 
          .B2(rModDataRead[7]), .B3(rModDataRead[6]), .CI(mco_15), .P0(mult_8u_9u_0_pp_3_15), 
          .P1(mult_8u_9u_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    AND2 AND2_t0_adj_214 (.A(SpriteRead_yInSprite[0]), .B(\currSprite_size[6] ), 
         .Z(mult_8u_8u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(125[10:63])
    AND2 AND2_t1_adj_215 (.A(SpriteRead_yInSprite[0]), .B(\currSprite_size[4] ), 
         .Z(mult_8u_8u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(123[10:63])
    AND2 AND2_t2_adj_216 (.A(SpriteRead_yInSprite[0]), .B(\currSprite_size[2] ), 
         .Z(mult_8u_8u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(121[10:63])
    AND2 AND2_t3_adj_217 (.A(SpriteRead_yInSprite[0]), .B(n17394), .Z(\Sprite_readAddr_13__N_752[0] )) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(119[10:63])
    FADD2B mult_8u_8u_0_Cadd_0_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(mult_8u_8u_0_pp_0_9)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_Cadd_2_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(mult_8u_8u_0_pp_1_11)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_Cadd_4_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(mult_8u_8u_0_pp_2_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B Cadd_mult_8u_8u_0_0_1 (.A0(GND_net), .A1(mult_8u_8u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_8u_8u_0_0_1), 
           .S1(\Sprite_readAddr_13__N_752[2] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_0_2 (.A0(mult_8u_8u_0_pp_0_3), .A1(mult_8u_8u_0_pp_0_4), 
           .B0(mult_8u_8u_0_pp_1_3), .B1(mult_8u_8u_0_pp_1_4), .CI(co_mult_8u_8u_0_0_1), 
           .COUT(co_mult_8u_8u_0_0_2), .S0(\Sprite_readAddr_13__N_752[3] ), 
           .S1(s_mult_8u_8u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_0_3 (.A0(mult_8u_8u_0_pp_0_5), .A1(mult_8u_8u_0_pp_0_6), 
           .B0(mult_8u_8u_0_pp_1_5), .B1(mult_8u_8u_0_pp_1_6), .CI(co_mult_8u_8u_0_0_2), 
           .COUT(co_mult_8u_8u_0_0_3), .S0(s_mult_8u_8u_0_0_5), .S1(s_mult_8u_8u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_0_4 (.A0(mult_8u_8u_0_pp_0_7), .A1(mult_8u_8u_0_pp_0_8), 
           .B0(mult_8u_8u_0_pp_1_7), .B1(mult_8u_8u_0_pp_1_8), .CI(co_mult_8u_8u_0_0_3), 
           .COUT(co_mult_8u_8u_0_0_4), .S0(s_mult_8u_8u_0_0_7), .S1(s_mult_8u_8u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_0_5 (.A0(mult_8u_8u_0_pp_0_9), .A1(GND_net), 
           .B0(mult_8u_8u_0_pp_1_9), .B1(mult_8u_8u_0_pp_1_10), .CI(co_mult_8u_8u_0_0_4), 
           .COUT(co_mult_8u_8u_0_0_5), .S0(s_mult_8u_8u_0_0_9), .S1(s_mult_8u_8u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_0_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_8u_0_pp_1_11), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_0_5), .COUT(co_mult_8u_8u_0_0_6), 
           .S0(s_mult_8u_8u_0_0_11), .S1(s_mult_8u_8u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B Cadd_mult_8u_8u_0_0_7 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_0_6), .S0(s_mult_8u_8u_0_0_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B Cadd_mult_8u_8u_0_1_1 (.A0(GND_net), .A1(mult_8u_8u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_8u_8u_0_1_1), 
           .S1(s_mult_8u_8u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_1_2 (.A0(mult_8u_8u_0_pp_2_7), .A1(mult_8u_8u_0_pp_2_8), 
           .B0(mult_8u_8u_0_pp_3_7), .B1(mult_8u_8u_0_pp_3_8), .CI(co_mult_8u_8u_0_1_1), 
           .COUT(co_mult_8u_8u_0_1_2), .S0(s_mult_8u_8u_0_1_7), .S1(s_mult_8u_8u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_1_3 (.A0(mult_8u_8u_0_pp_2_9), .A1(mult_8u_8u_0_pp_2_10), 
           .B0(mult_8u_8u_0_pp_3_9), .B1(mult_8u_8u_0_pp_3_10), .CI(co_mult_8u_8u_0_1_2), 
           .COUT(co_mult_8u_8u_0_1_3), .S0(s_mult_8u_8u_0_1_9), .S1(s_mult_8u_8u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_1_4 (.A0(mult_8u_8u_0_pp_2_11), .A1(mult_8u_8u_0_pp_2_12), 
           .B0(mult_8u_8u_0_pp_3_11), .B1(mult_8u_8u_0_pp_3_12), .CI(co_mult_8u_8u_0_1_3), 
           .COUT(co_mult_8u_8u_0_1_4), .S0(s_mult_8u_8u_0_1_11), .S1(s_mult_8u_8u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B mult_8u_8u_0_add_1_5 (.A0(mult_8u_8u_0_pp_2_13), .A1(GND_net), 
           .B0(mult_8u_8u_0_pp_3_13), .B1(mult_8u_8u_0_pp_3_14), .CI(co_mult_8u_8u_0_1_4), 
           .S0(s_mult_8u_8u_0_1_13), .S1(s_mult_8u_8u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B Cadd_t_mult_8u_8u_0_2_1 (.A0(GND_net), .A1(s_mult_8u_8u_0_0_4), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_2_4), .CI(GND_net), .COUT(co_t_mult_8u_8u_0_2_1), 
           .S1(\Sprite_readAddr_13__N_752[4] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B t_mult_8u_8u_0_add_2_2 (.A0(s_mult_8u_8u_0_0_5), .A1(s_mult_8u_8u_0_0_6), 
           .B0(mult_8u_8u_0_pp_2_5), .B1(s_mult_8u_8u_0_1_6), .CI(co_t_mult_8u_8u_0_2_1), 
           .COUT(co_t_mult_8u_8u_0_2_2), .S0(\Sprite_readAddr_13__N_752[5] ), 
           .S1(\Sprite_readAddr_13__N_752[6] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B t_mult_8u_8u_0_add_2_3 (.A0(s_mult_8u_8u_0_0_7), .A1(s_mult_8u_8u_0_0_8), 
           .B0(s_mult_8u_8u_0_1_7), .B1(s_mult_8u_8u_0_1_8), .CI(co_t_mult_8u_8u_0_2_2), 
           .COUT(co_t_mult_8u_8u_0_2_3), .S0(\Sprite_readAddr_13__N_752[7] ), 
           .S1(\Sprite_readAddr_13__N_752[8] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B t_mult_8u_8u_0_add_2_4 (.A0(s_mult_8u_8u_0_0_9), .A1(s_mult_8u_8u_0_0_10), 
           .B0(s_mult_8u_8u_0_1_9), .B1(s_mult_8u_8u_0_1_10), .CI(co_t_mult_8u_8u_0_2_3), 
           .COUT(co_t_mult_8u_8u_0_2_4), .S0(\Sprite_readAddr_13__N_752[9] ), 
           .S1(\Sprite_readAddr_13__N_752[10] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B t_mult_8u_8u_0_add_2_5 (.A0(s_mult_8u_8u_0_0_11), .A1(s_mult_8u_8u_0_0_12), 
           .B0(s_mult_8u_8u_0_1_11), .B1(s_mult_8u_8u_0_1_12), .CI(co_t_mult_8u_8u_0_2_4), 
           .COUT(co_t_mult_8u_8u_0_2_5), .S0(\Sprite_readAddr_13__N_752[11] ), 
           .S1(\Sprite_readAddr_13__N_752[12] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    FADD2B t_mult_8u_8u_0_add_2_6 (.A0(s_mult_8u_8u_0_0_13), .A1(GND_net), 
           .B0(s_mult_8u_8u_0_1_13), .B1(s_mult_8u_8u_0_1_14), .CI(co_t_mult_8u_8u_0_2_5), 
           .S0(\Sprite_readAddr_13__N_752[13] )) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_0_0 (.A0(SpriteRead_yInSprite[0]), .A1(SpriteRead_yInSprite[1]), 
          .A2(SpriteRead_yInSprite[1]), .A3(SpriteRead_yInSprite[2]), .B0(\currSprite_size[1] ), 
          .B1(n17394), .B2(\currSprite_size[1] ), .B3(n17394), .CI(mult_8u_8u_0_cin_lr_0), 
          .CO(mco_adj_1775), .P0(\Sprite_readAddr_13__N_752[1] ), .P1(mult_8u_8u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_0_1 (.A0(SpriteRead_yInSprite[2]), .A1(SpriteRead_yInSprite[3]), 
          .A2(SpriteRead_yInSprite[3]), .A3(SpriteRead_yInSprite[4]), .B0(\currSprite_size[1] ), 
          .B1(n17394), .B2(\currSprite_size[1] ), .B3(n17394), .CI(mco_adj_1775), 
          .CO(mco_1_adj_1776), .P0(mult_8u_8u_0_pp_0_3), .P1(mult_8u_8u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_0_2 (.A0(SpriteRead_yInSprite[4]), .A1(SpriteRead_yInSprite[5]), 
          .A2(SpriteRead_yInSprite[5]), .A3(SpriteRead_yInSprite[6]), .B0(\currSprite_size[1] ), 
          .B1(n17394), .B2(\currSprite_size[1] ), .B3(n17394), .CI(mco_1_adj_1776), 
          .CO(mco_2_adj_1777), .P0(mult_8u_8u_0_pp_0_5), .P1(mult_8u_8u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_0_3 (.A0(SpriteRead_yInSprite[6]), .A1(SpriteRead_yInSprite[7]), 
          .A2(SpriteRead_yInSprite[7]), .A3(GND_net), .B0(\currSprite_size[1] ), 
          .B1(n17394), .B2(\currSprite_size[1] ), .B3(n17394), .CI(mco_2_adj_1777), 
          .CO(mfco), .P0(mult_8u_8u_0_pp_0_7), .P1(mult_8u_8u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_2_0 (.A0(SpriteRead_yInSprite[0]), .A1(SpriteRead_yInSprite[1]), 
          .A2(SpriteRead_yInSprite[1]), .A3(SpriteRead_yInSprite[2]), .B0(\currSprite_size[3] ), 
          .B1(\currSprite_size[2] ), .B2(\currSprite_size[3] ), .B3(\currSprite_size[2] ), 
          .CI(mult_8u_8u_0_cin_lr_2), .CO(mco_3_adj_1778), .P0(mult_8u_8u_0_pp_1_3), 
          .P1(mult_8u_8u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_2_1 (.A0(SpriteRead_yInSprite[2]), .A1(SpriteRead_yInSprite[3]), 
          .A2(SpriteRead_yInSprite[3]), .A3(SpriteRead_yInSprite[4]), .B0(\currSprite_size[3] ), 
          .B1(\currSprite_size[2] ), .B2(\currSprite_size[3] ), .B3(\currSprite_size[2] ), 
          .CI(mco_3_adj_1778), .CO(mco_4_adj_1779), .P0(mult_8u_8u_0_pp_1_5), 
          .P1(mult_8u_8u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_2_2 (.A0(SpriteRead_yInSprite[4]), .A1(SpriteRead_yInSprite[5]), 
          .A2(SpriteRead_yInSprite[5]), .A3(SpriteRead_yInSprite[6]), .B0(\currSprite_size[3] ), 
          .B1(\currSprite_size[2] ), .B2(\currSprite_size[3] ), .B3(\currSprite_size[2] ), 
          .CI(mco_4_adj_1779), .CO(mco_5_adj_1780), .P0(mult_8u_8u_0_pp_1_7), 
          .P1(mult_8u_8u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_2_3 (.A0(SpriteRead_yInSprite[6]), .A1(SpriteRead_yInSprite[7]), 
          .A2(SpriteRead_yInSprite[7]), .A3(GND_net), .B0(\currSprite_size[3] ), 
          .B1(\currSprite_size[2] ), .B2(\currSprite_size[3] ), .B3(\currSprite_size[2] ), 
          .CI(mco_5_adj_1780), .CO(mfco_1), .P0(mult_8u_8u_0_pp_1_9), 
          .P1(mult_8u_8u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_4_0 (.A0(SpriteRead_yInSprite[0]), .A1(SpriteRead_yInSprite[1]), 
          .A2(SpriteRead_yInSprite[1]), .A3(SpriteRead_yInSprite[2]), .B0(\currSprite_size[5] ), 
          .B1(\currSprite_size[4] ), .B2(\currSprite_size[5] ), .B3(\currSprite_size[4] ), 
          .CI(mult_8u_8u_0_cin_lr_4), .CO(mco_6_adj_1781), .P0(mult_8u_8u_0_pp_2_5), 
          .P1(mult_8u_8u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_4_1 (.A0(SpriteRead_yInSprite[2]), .A1(SpriteRead_yInSprite[3]), 
          .A2(SpriteRead_yInSprite[3]), .A3(SpriteRead_yInSprite[4]), .B0(\currSprite_size[5] ), 
          .B1(\currSprite_size[4] ), .B2(\currSprite_size[5] ), .B3(\currSprite_size[4] ), 
          .CI(mco_6_adj_1781), .CO(mco_7_adj_1782), .P0(mult_8u_8u_0_pp_2_7), 
          .P1(mult_8u_8u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_4_2 (.A0(SpriteRead_yInSprite[4]), .A1(SpriteRead_yInSprite[5]), 
          .A2(SpriteRead_yInSprite[5]), .A3(SpriteRead_yInSprite[6]), .B0(\currSprite_size[5] ), 
          .B1(\currSprite_size[4] ), .B2(\currSprite_size[5] ), .B3(\currSprite_size[4] ), 
          .CI(mco_7_adj_1782), .CO(mco_8_adj_1783), .P0(mult_8u_8u_0_pp_2_9), 
          .P1(mult_8u_8u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_4_3 (.A0(SpriteRead_yInSprite[6]), .A1(SpriteRead_yInSprite[7]), 
          .A2(SpriteRead_yInSprite[7]), .A3(GND_net), .B0(\currSprite_size[5] ), 
          .B1(\currSprite_size[4] ), .B2(\currSprite_size[5] ), .B3(\currSprite_size[4] ), 
          .CI(mco_8_adj_1783), .CO(mfco_2), .P0(mult_8u_8u_0_pp_2_11), 
          .P1(mult_8u_8u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_6_0 (.A0(SpriteRead_yInSprite[0]), .A1(SpriteRead_yInSprite[1]), 
          .A2(SpriteRead_yInSprite[1]), .A3(SpriteRead_yInSprite[2]), .B0(\currSprite_size[7] ), 
          .B1(\currSprite_size[6] ), .B2(\currSprite_size[7] ), .B3(\currSprite_size[6] ), 
          .CI(mult_8u_8u_0_cin_lr_6), .CO(mco_9_adj_1784), .P0(mult_8u_8u_0_pp_3_7), 
          .P1(mult_8u_8u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_6_1 (.A0(SpriteRead_yInSprite[2]), .A1(SpriteRead_yInSprite[3]), 
          .A2(SpriteRead_yInSprite[3]), .A3(SpriteRead_yInSprite[4]), .B0(\currSprite_size[7] ), 
          .B1(\currSprite_size[6] ), .B2(\currSprite_size[7] ), .B3(\currSprite_size[6] ), 
          .CI(mco_9_adj_1784), .CO(mco_10_adj_1785), .P0(mult_8u_8u_0_pp_3_9), 
          .P1(mult_8u_8u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_6_2 (.A0(SpriteRead_yInSprite[4]), .A1(SpriteRead_yInSprite[5]), 
          .A2(SpriteRead_yInSprite[5]), .A3(SpriteRead_yInSprite[6]), .B0(\currSprite_size[7] ), 
          .B1(\currSprite_size[6] ), .B2(\currSprite_size[7] ), .B3(\currSprite_size[6] ), 
          .CI(mco_10_adj_1785), .CO(mco_11_adj_1786), .P0(mult_8u_8u_0_pp_3_11), 
          .P1(mult_8u_8u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    MULT2 mult_8u_8u_0_mult_6_3 (.A0(SpriteRead_yInSprite[6]), .A1(SpriteRead_yInSprite[7]), 
          .A2(SpriteRead_yInSprite[7]), .A3(GND_net), .B0(\currSprite_size[7] ), 
          .B1(\currSprite_size[6] ), .B2(\currSprite_size[7] ), .B3(\currSprite_size[6] ), 
          .CI(mco_11_adj_1786), .P0(mult_8u_8u_0_pp_3_13), .P1(mult_8u_8u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(274[71:97])
    CCU2D add_319_9 (.A0(rModDataTrans[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14117), .S0(rModDataWrite_15__N_1670[7]), .S1(rModDataWrite_15__N_1670[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_319_9.INIT0 = 16'hf555;
    defparam add_319_9.INIT1 = 16'h0000;
    defparam add_319_9.INJECT1_0 = "NO";
    defparam add_319_9.INJECT1_1 = "NO";
    CCU2D add_319_7 (.A0(rModDataTrans[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(rModDataTrans[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14116), .COUT(n14117), .S0(rModDataWrite_15__N_1670[5]), 
          .S1(rModDataWrite_15__N_1670[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_319_7.INIT0 = 16'hf555;
    defparam add_319_7.INIT1 = 16'hf555;
    defparam add_319_7.INJECT1_0 = "NO";
    defparam add_319_7.INJECT1_1 = "NO";
    CCU2D add_319_5 (.A0(rModDataTrans[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(rModDataTrans[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14115), .COUT(n14116), .S0(rModDataWrite_15__N_1670[3]), 
          .S1(rModDataWrite_15__N_1670[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_319_5.INIT0 = 16'hf555;
    defparam add_319_5.INIT1 = 16'hf555;
    defparam add_319_5.INJECT1_0 = "NO";
    defparam add_319_5.INJECT1_1 = "NO";
    CCU2D add_319_3 (.A0(rModDataTrans[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(rModDataTrans[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14114), .COUT(n14115), .S0(rModDataWrite_15__N_1670[1]), 
          .S1(rModDataWrite_15__N_1670[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_319_3.INIT0 = 16'hf555;
    defparam add_319_3.INIT1 = 16'hf555;
    defparam add_319_3.INJECT1_0 = "NO";
    defparam add_319_3.INJECT1_1 = "NO";
    AND2 AND2_t0_adj_218 (.A(data[0]), .B(rModDataTrans[6]), .Z(mult_8u_8u_0_pp_3_6_adj_1787)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(125[10:63])
    AND2 AND2_t1_adj_219 (.A(data[0]), .B(rModDataTrans[4]), .Z(mult_8u_8u_0_pp_2_4_adj_1788)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(123[10:63])
    AND2 AND2_t2_adj_220 (.A(data[0]), .B(rModDataTrans[2]), .Z(mult_8u_8u_0_pp_1_2_adj_1789)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(121[10:63])
    AND2 AND2_t3_adj_221 (.A(data[0]), .B(rModDataTrans[0]), .Z(rModDataWrite_15__N_1637[0])) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(119[10:63])
    FADD2B mult_8u_8u_0_Cadd_0_4_adj_222 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_adj_1791), .S0(mult_8u_8u_0_pp_0_9_adj_1790)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_cin_lr_add_2_adj_223 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_2_adj_1792)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_Cadd_2_4_adj_224 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1_adj_1794), .S0(mult_8u_8u_0_pp_1_11_adj_1793)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_cin_lr_add_4_adj_225 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_4_adj_1795)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_Cadd_4_4_adj_226 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2_adj_1797), .S0(mult_8u_8u_0_pp_2_13_adj_1796)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_cin_lr_add_6_adj_227 (.A0(GND_net), .A1(GND_net), 
           .B0(GND_net), .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_6_adj_1798)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_Cadd_6_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(mult_8u_8u_0_pp_3_15)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_mult_8u_8u_0_0_1_adj_228 (.A0(GND_net), .A1(mult_8u_8u_0_pp_0_2_adj_1800), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_1_2_adj_1789), .CI(GND_net), 
           .COUT(co_mult_8u_8u_0_0_1_adj_1799), .S1(rModDataWrite_15__N_1637[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_2_adj_229 (.A0(mult_8u_8u_0_pp_0_3_adj_1804), 
           .A1(mult_8u_8u_0_pp_0_4_adj_1803), .B0(mult_8u_8u_0_pp_1_3_adj_1806), 
           .B1(mult_8u_8u_0_pp_1_4_adj_1805), .CI(co_mult_8u_8u_0_0_1_adj_1799), 
           .COUT(co_mult_8u_8u_0_0_2_adj_1801), .S0(rModDataWrite_15__N_1637[3]), 
           .S1(s_mult_8u_8u_0_0_4_adj_1802)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_3_adj_230 (.A0(mult_8u_8u_0_pp_0_5_adj_1811), 
           .A1(mult_8u_8u_0_pp_0_6_adj_1810), .B0(mult_8u_8u_0_pp_1_5_adj_1813), 
           .B1(mult_8u_8u_0_pp_1_6_adj_1812), .CI(co_mult_8u_8u_0_0_2_adj_1801), 
           .COUT(co_mult_8u_8u_0_0_3_adj_1807), .S0(s_mult_8u_8u_0_0_5_adj_1808), 
           .S1(s_mult_8u_8u_0_0_6_adj_1809)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_4_adj_231 (.A0(mult_8u_8u_0_pp_0_7_adj_1818), 
           .A1(mult_8u_8u_0_pp_0_8_adj_1817), .B0(mult_8u_8u_0_pp_1_7_adj_1820), 
           .B1(mult_8u_8u_0_pp_1_8_adj_1819), .CI(co_mult_8u_8u_0_0_3_adj_1807), 
           .COUT(co_mult_8u_8u_0_0_4_adj_1814), .S0(s_mult_8u_8u_0_0_7_adj_1815), 
           .S1(s_mult_8u_8u_0_0_8_adj_1816)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_5_adj_232 (.A0(mult_8u_8u_0_pp_0_9_adj_1790), 
           .A1(GND_net), .B0(mult_8u_8u_0_pp_1_9_adj_1825), .B1(mult_8u_8u_0_pp_1_10_adj_1824), 
           .CI(co_mult_8u_8u_0_0_4_adj_1814), .COUT(co_mult_8u_8u_0_0_5_adj_1821), 
           .S0(s_mult_8u_8u_0_0_9_adj_1822), .S1(s_mult_8u_8u_0_0_10_adj_1823)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_6_adj_233 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_8u_0_pp_1_11_adj_1793), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_0_5_adj_1821), .COUT(co_mult_8u_8u_0_0_6_adj_1826), 
           .S0(s_mult_8u_8u_0_0_11_adj_1827), .S1(s_mult_8u_8u_0_0_12_adj_1828)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_mult_8u_8u_0_0_7_adj_234 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_0_6_adj_1826), .S0(s_mult_8u_8u_0_0_13_adj_1829)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_mult_8u_8u_0_1_1_adj_235 (.A0(GND_net), .A1(mult_8u_8u_0_pp_2_6_adj_1832), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_3_6_adj_1787), .CI(GND_net), 
           .COUT(co_mult_8u_8u_0_1_1_adj_1830), .S1(s_mult_8u_8u_0_1_6_adj_1831)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_2_adj_236 (.A0(mult_8u_8u_0_pp_2_7_adj_1837), 
           .A1(mult_8u_8u_0_pp_2_8_adj_1836), .B0(mult_8u_8u_0_pp_3_7_adj_1839), 
           .B1(mult_8u_8u_0_pp_3_8_adj_1838), .CI(co_mult_8u_8u_0_1_1_adj_1830), 
           .COUT(co_mult_8u_8u_0_1_2_adj_1833), .S0(s_mult_8u_8u_0_1_7_adj_1834), 
           .S1(s_mult_8u_8u_0_1_8_adj_1835)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_3_adj_237 (.A0(mult_8u_8u_0_pp_2_9_adj_1844), 
           .A1(mult_8u_8u_0_pp_2_10_adj_1843), .B0(mult_8u_8u_0_pp_3_9_adj_1846), 
           .B1(mult_8u_8u_0_pp_3_10_adj_1845), .CI(co_mult_8u_8u_0_1_2_adj_1833), 
           .COUT(co_mult_8u_8u_0_1_3_adj_1840), .S0(s_mult_8u_8u_0_1_9_adj_1841), 
           .S1(s_mult_8u_8u_0_1_10_adj_1842)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_4_adj_238 (.A0(mult_8u_8u_0_pp_2_11_adj_1851), 
           .A1(mult_8u_8u_0_pp_2_12_adj_1850), .B0(mult_8u_8u_0_pp_3_11_adj_1853), 
           .B1(mult_8u_8u_0_pp_3_12_adj_1852), .CI(co_mult_8u_8u_0_1_3_adj_1840), 
           .COUT(co_mult_8u_8u_0_1_4_adj_1847), .S0(s_mult_8u_8u_0_1_11_adj_1848), 
           .S1(s_mult_8u_8u_0_1_12_adj_1849)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_5_adj_239 (.A0(mult_8u_8u_0_pp_2_13_adj_1796), 
           .A1(GND_net), .B0(mult_8u_8u_0_pp_3_13_adj_1857), .B1(mult_8u_8u_0_pp_3_14_adj_1856), 
           .CI(co_mult_8u_8u_0_1_4_adj_1847), .COUT(co_mult_8u_8u_0_1_5), 
           .S0(s_mult_8u_8u_0_1_13_adj_1854), .S1(s_mult_8u_8u_0_1_14_adj_1855)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_8u_0_pp_3_15), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_1_5), .S0(s_mult_8u_8u_0_1_15)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_t_mult_8u_8u_0_2_1_adj_240 (.A0(GND_net), .A1(s_mult_8u_8u_0_0_4_adj_1802), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_2_4_adj_1788), .CI(GND_net), 
           .COUT(co_t_mult_8u_8u_0_2_1_adj_1858), .S1(rModDataWrite_15__N_1637[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_2_adj_241 (.A0(s_mult_8u_8u_0_0_5_adj_1808), 
           .A1(s_mult_8u_8u_0_0_6_adj_1809), .B0(mult_8u_8u_0_pp_2_5_adj_1860), 
           .B1(s_mult_8u_8u_0_1_6_adj_1831), .CI(co_t_mult_8u_8u_0_2_1_adj_1858), 
           .COUT(co_t_mult_8u_8u_0_2_2_adj_1859), .S0(rModDataWrite_15__N_1637[5]), 
           .S1(rModDataWrite_15__N_1637[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_3_adj_242 (.A0(s_mult_8u_8u_0_0_7_adj_1815), 
           .A1(s_mult_8u_8u_0_0_8_adj_1816), .B0(s_mult_8u_8u_0_1_7_adj_1834), 
           .B1(s_mult_8u_8u_0_1_8_adj_1835), .CI(co_t_mult_8u_8u_0_2_2_adj_1859), 
           .COUT(co_t_mult_8u_8u_0_2_3_adj_1861), .S0(rModDataWrite_15__N_1637[7]), 
           .S1(rModDataWrite_15__N_1637[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_4_adj_243 (.A0(s_mult_8u_8u_0_0_9_adj_1822), 
           .A1(s_mult_8u_8u_0_0_10_adj_1823), .B0(s_mult_8u_8u_0_1_9_adj_1841), 
           .B1(s_mult_8u_8u_0_1_10_adj_1842), .CI(co_t_mult_8u_8u_0_2_3_adj_1861), 
           .COUT(co_t_mult_8u_8u_0_2_4_adj_1862), .S0(rModDataWrite_15__N_1637[9]), 
           .S1(rModDataWrite_15__N_1637[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_5_adj_244 (.A0(s_mult_8u_8u_0_0_11_adj_1827), 
           .A1(s_mult_8u_8u_0_0_12_adj_1828), .B0(s_mult_8u_8u_0_1_11_adj_1848), 
           .B1(s_mult_8u_8u_0_1_12_adj_1849), .CI(co_t_mult_8u_8u_0_2_4_adj_1862), 
           .COUT(co_t_mult_8u_8u_0_2_5_adj_1863), .S0(rModDataWrite_15__N_1637[11]), 
           .S1(rModDataWrite_15__N_1637[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_6_adj_245 (.A0(s_mult_8u_8u_0_0_13_adj_1829), 
           .A1(GND_net), .B0(s_mult_8u_8u_0_1_13_adj_1854), .B1(s_mult_8u_8u_0_1_14_adj_1855), 
           .CI(co_t_mult_8u_8u_0_2_5_adj_1863), .COUT(co_t_mult_8u_8u_0_2_6), 
           .S0(rModDataWrite_15__N_1637[13]), .S1(rModDataWrite_15__N_1637[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_7 (.A0(GND_net), .A1(GND_net), .B0(s_mult_8u_8u_0_1_15), 
           .B1(GND_net), .CI(co_t_mult_8u_8u_0_2_6), .S0(rModDataWrite_15__N_1637[15])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_0_adj_246 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mult_8u_8u_0_cin_lr_0_adj_1773), 
          .CO(mco_adj_1864), .P0(rModDataWrite_15__N_1637[1]), .P1(mult_8u_8u_0_pp_0_2_adj_1800)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_1_adj_247 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mco_adj_1864), 
          .CO(mco_1_adj_1865), .P0(mult_8u_8u_0_pp_0_3_adj_1804), .P1(mult_8u_8u_0_pp_0_4_adj_1803)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_2_adj_248 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mco_1_adj_1865), 
          .CO(mco_2_adj_1866), .P0(mult_8u_8u_0_pp_0_5_adj_1811), .P1(mult_8u_8u_0_pp_0_6_adj_1810)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_3_adj_249 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mco_2_adj_1866), 
          .CO(mfco_adj_1791), .P0(mult_8u_8u_0_pp_0_7_adj_1818), .P1(mult_8u_8u_0_pp_0_8_adj_1817)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_0_adj_250 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mult_8u_8u_0_cin_lr_2_adj_1792), 
          .CO(mco_3_adj_1867), .P0(mult_8u_8u_0_pp_1_3_adj_1806), .P1(mult_8u_8u_0_pp_1_4_adj_1805)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_1_adj_251 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mco_3_adj_1867), 
          .CO(mco_4_adj_1868), .P0(mult_8u_8u_0_pp_1_5_adj_1813), .P1(mult_8u_8u_0_pp_1_6_adj_1812)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_2_adj_252 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mco_4_adj_1868), 
          .CO(mco_5_adj_1869), .P0(mult_8u_8u_0_pp_1_7_adj_1820), .P1(mult_8u_8u_0_pp_1_8_adj_1819)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_3_adj_253 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mco_5_adj_1869), 
          .CO(mfco_1_adj_1794), .P0(mult_8u_8u_0_pp_1_9_adj_1825), .P1(mult_8u_8u_0_pp_1_10_adj_1824)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_0_adj_254 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mult_8u_8u_0_cin_lr_4_adj_1795), 
          .CO(mco_6_adj_1870), .P0(mult_8u_8u_0_pp_2_5_adj_1860), .P1(mult_8u_8u_0_pp_2_6_adj_1832)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_1_adj_255 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mco_6_adj_1870), 
          .CO(mco_7_adj_1871), .P0(mult_8u_8u_0_pp_2_7_adj_1837), .P1(mult_8u_8u_0_pp_2_8_adj_1836)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_2_adj_256 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mco_7_adj_1871), 
          .CO(mco_8_adj_1872), .P0(mult_8u_8u_0_pp_2_9_adj_1844), .P1(mult_8u_8u_0_pp_2_10_adj_1843)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_3_adj_257 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mco_8_adj_1872), 
          .CO(mfco_2_adj_1797), .P0(mult_8u_8u_0_pp_2_11_adj_1851), .P1(mult_8u_8u_0_pp_2_12_adj_1850)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_0_adj_258 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mult_8u_8u_0_cin_lr_6_adj_1798), 
          .CO(mco_9_adj_1873), .P0(mult_8u_8u_0_pp_3_7_adj_1839), .P1(mult_8u_8u_0_pp_3_8_adj_1838)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_1_adj_259 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mco_9_adj_1873), 
          .CO(mco_10_adj_1874), .P0(mult_8u_8u_0_pp_3_9_adj_1846), .P1(mult_8u_8u_0_pp_3_10_adj_1845)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_2_adj_260 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mco_10_adj_1874), 
          .CO(mco_11_adj_1875), .P0(mult_8u_8u_0_pp_3_11_adj_1853), .P1(mult_8u_8u_0_pp_3_12_adj_1852)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_3_adj_261 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mco_11_adj_1875), 
          .CO(mfco_3), .P0(mult_8u_8u_0_pp_3_13_adj_1857), .P1(mult_8u_8u_0_pp_3_14_adj_1856)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    CCU2D add_319_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(rModDataTrans[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n14114), .S1(rModDataWrite_15__N_1670[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_319_1.INIT0 = 16'hF000;
    defparam add_319_1.INIT1 = 16'h0aaa;
    defparam add_319_1.INJECT1_0 = "NO";
    defparam add_319_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_262 (.A(n9_adj_1876), .B(n17270), .C(n14_adj_1877), 
         .D(n10_adj_1878), .Z(LOGIC_CLOCK_enable_80)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_4_lut_adj_262.init = 16'h8000;
    LUT4 i1_2_lut (.A(state_c[3]), .B(state_c[6]), .Z(n9_adj_1876)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_263 (.A(state[1]), .B(state_c[7]), .C(state[4]), 
         .D(state_c[2]), .Z(n14_adj_1877)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i6_4_lut_adj_263.init = 16'h8000;
    LUT4 i2_2_lut_adj_264 (.A(state_c[5]), .B(state_c[0]), .Z(n10_adj_1878)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i2_2_lut_adj_264.init = 16'h8888;
    FD1P3AX transferMode_i0_i1 (.D(\BUS_data[1] ), .SP(LOGIC_CLOCK_enable_216), 
            .CK(LOGIC_CLOCK), .Q(transferMode[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i1.GSR = "DISABLED";
    FD1P3AX transferMode_i0_i2 (.D(\BUS_data[2] ), .SP(LOGIC_CLOCK_enable_216), 
            .CK(LOGIC_CLOCK), .Q(transferMode[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i2.GSR = "DISABLED";
    FD1P3AX transferMode_i0_i3 (.D(\BUS_data[3] ), .SP(LOGIC_CLOCK_enable_216), 
            .CK(LOGIC_CLOCK), .Q(transferMode[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i3.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i2 (.D(PIC_ADDR_IN_c_1), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i2.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i3 (.D(PIC_ADDR_IN_c_2), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i3.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i4 (.D(PIC_ADDR_IN_c_3), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i4.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i5 (.D(PIC_ADDR_IN_c_4), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i5.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i6 (.D(PIC_ADDR_IN_c_5), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i6.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i7 (.D(PIC_ADDR_IN_c_6), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i7.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i8 (.D(PIC_ADDR_IN_c_7), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i8.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i9 (.D(PIC_ADDR_IN_c_8), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i9.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i10 (.D(PIC_ADDR_IN_c_9), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i10.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i11 (.D(PIC_ADDR_IN_c_10), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i11.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i12 (.D(PIC_ADDR_IN_c_11), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i12.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i13 (.D(PIC_ADDR_IN_c_12), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i13.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i14 (.D(PIC_ADDR_IN_c_13), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i14.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i15 (.D(PIC_ADDR_IN_c_14), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i15.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i16 (.D(PIC_ADDR_IN_c_15), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i16.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i17 (.D(PIC_ADDR_IN_c_16), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i17.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i18 (.D(PIC_ADDR_IN_c_17), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i18.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i19 (.D(PIC_ADDR_IN_c_18), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i19.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i1 (.D(\BUS_data[1] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i1.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i2 (.D(\BUS_data[2] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i2.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i3 (.D(\BUS_data[3] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i3.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i4 (.D(\BUS_data[4] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i4.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i5 (.D(\BUS_data[5] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i5.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i6 (.D(\BUS_data[6] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i6.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i7 (.D(\BUS_data[7] ), .SP(LOGIC_CLOCK_enable_241), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i7.GSR = "DISABLED";
    FD1P3AX writeData_i0_i1 (.D(writeData_15__N_1719[1]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(writeData_c[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i1.GSR = "DISABLED";
    FD1P3AX writeData_i0_i2 (.D(writeData_15__N_1719[2]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(writeData_c[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i2.GSR = "DISABLED";
    FD1P3AX writeData_i0_i3 (.D(writeData_15__N_1719[3]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(writeData_c[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i3.GSR = "DISABLED";
    FD1P3AX writeData_i0_i4 (.D(writeData_15__N_1719[4]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(\writeData[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i4.GSR = "DISABLED";
    FD1P3AX writeData_i0_i5 (.D(writeData_15__N_1719[5]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(\writeData[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i5.GSR = "DISABLED";
    FD1P3AX writeData_i0_i6 (.D(writeData_15__N_1719[6]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(\writeData[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i6.GSR = "DISABLED";
    FD1P3AX writeData_i0_i7 (.D(writeData_15__N_1719[7]), .SP(LOGIC_CLOCK_enable_248), 
            .CK(LOGIC_CLOCK), .Q(\writeData[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i7.GSR = "DISABLED";
    FD1S3DX state_i1 (.D(state_7__N_1600[1]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_1547), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i1.GSR = "DISABLED";
    FD1P3DX state_i2 (.D(n18280), .SP(LOGIC_CLOCK_enable_249), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_1547), .Q(state_c[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i2.GSR = "DISABLED";
    FD1P3DX state_i3 (.D(n18280), .SP(LOGIC_CLOCK_enable_250), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_1547), .Q(state_c[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i3.GSR = "DISABLED";
    FD1S3DX state_i4 (.D(state_7__N_1600[4]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_1547), 
            .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i4.GSR = "DISABLED";
    FD1P3DX state_i5 (.D(n18280), .SP(LOGIC_CLOCK_enable_251), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_1547), .Q(state_c[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i5.GSR = "DISABLED";
    FD1P3DX state_i6 (.D(n18280), .SP(LOGIC_CLOCK_enable_252), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_1547), .Q(state_c[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i6.GSR = "DISABLED";
    FD1S3DX state_i7 (.D(state_7__N_1600[7]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_1547), 
            .Q(state_c[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i7.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i1 (.D(data[9]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i1.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i2 (.D(data[10]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i2.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i3 (.D(data[11]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i3.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i4 (.D(data[12]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i4.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i5 (.D(data[13]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i5.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i6 (.D(data[14]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i6.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i7 (.D(data[15]), .SP(LOGIC_CLOCK_enable_259), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=218, LSE_RLINE=218 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i7.GSR = "DISABLED";
    CCU2D add_320_16 (.A0(rModDataWrite_15__N_1620[14]), .B0(rModDataWrite_15__N_1637[14]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[15]), 
          .B1(rModDataWrite_15__N_1637[15]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14103), .S0(rModDataWrite[14]), .S1(rModDataWrite[15]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_16.INIT0 = 16'h5666;
    defparam add_320_16.INIT1 = 16'h5666;
    defparam add_320_16.INJECT1_0 = "NO";
    defparam add_320_16.INJECT1_1 = "NO";
    LUT4 i6620_2_lut (.A(PIC_DATA_IN_out_0), .B(PIC_WE_IN_c), .Z(data[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6620_2_lut.init = 16'h2222;
    LUT4 i6868_2_lut (.A(PIC_DATA_IN_out_2), .B(PIC_WE_IN_c), .Z(data[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6868_2_lut.init = 16'h2222;
    CCU2D add_320_14 (.A0(rModDataWrite_15__N_1620[12]), .B0(rModDataWrite_15__N_1637[12]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[13]), 
          .B1(rModDataWrite_15__N_1637[13]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14102), .COUT(n14103), .S0(rModDataWrite[12]), .S1(rModDataWrite[13]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_14.INIT0 = 16'h5666;
    defparam add_320_14.INIT1 = 16'h5666;
    defparam add_320_14.INJECT1_0 = "NO";
    defparam add_320_14.INJECT1_1 = "NO";
    CCU2D add_320_12 (.A0(rModDataWrite_15__N_1620[10]), .B0(rModDataWrite_15__N_1637[10]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[11]), 
          .B1(rModDataWrite_15__N_1637[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14101), .COUT(n14102), .S0(rModDataWrite[10]), .S1(rModDataWrite[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_12.INIT0 = 16'h5666;
    defparam add_320_12.INIT1 = 16'h5666;
    defparam add_320_12.INJECT1_0 = "NO";
    defparam add_320_12.INJECT1_1 = "NO";
    CCU2D add_320_10 (.A0(rModDataWrite_15__N_1620[8]), .B0(rModDataWrite_15__N_1637[8]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[9]), 
          .B1(rModDataWrite_15__N_1637[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14100), .COUT(n14101), .S0(rModDataWrite[8]), .S1(rModDataWrite[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_10.INIT0 = 16'h5666;
    defparam add_320_10.INIT1 = 16'h5666;
    defparam add_320_10.INJECT1_0 = "NO";
    defparam add_320_10.INJECT1_1 = "NO";
    LUT4 i6867_2_lut (.A(PIC_DATA_IN_out_1), .B(PIC_WE_IN_c), .Z(data[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6867_2_lut.init = 16'h2222;
    LUT4 i6870_2_lut (.A(PIC_DATA_IN_out_4), .B(PIC_WE_IN_c), .Z(data[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6870_2_lut.init = 16'h2222;
    LUT4 i6869_2_lut (.A(PIC_DATA_IN_out_3), .B(PIC_WE_IN_c), .Z(data[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6869_2_lut.init = 16'h2222;
    LUT4 i6872_2_lut (.A(PIC_DATA_IN_out_6), .B(PIC_WE_IN_c), .Z(data[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6872_2_lut.init = 16'h2222;
    CCU2D add_320_8 (.A0(rModDataWrite_15__N_1620[6]), .B0(rModDataWrite_15__N_1637[6]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[7]), 
          .B1(rModDataWrite_15__N_1637[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14099), .COUT(n14100));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_8.INIT0 = 16'h5666;
    defparam add_320_8.INIT1 = 16'h5666;
    defparam add_320_8.INJECT1_0 = "NO";
    defparam add_320_8.INJECT1_1 = "NO";
    LUT4 i6871_2_lut (.A(PIC_DATA_IN_out_5), .B(PIC_WE_IN_c), .Z(data[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6871_2_lut.init = 16'h2222;
    CCU2D add_320_6 (.A0(rModDataWrite_15__N_1620[4]), .B0(rModDataWrite_15__N_1637[4]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[5]), 
          .B1(rModDataWrite_15__N_1637[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14098), .COUT(n14099));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_6.INIT0 = 16'h5666;
    defparam add_320_6.INIT1 = 16'h5666;
    defparam add_320_6.INJECT1_0 = "NO";
    defparam add_320_6.INJECT1_1 = "NO";
    CCU2D add_320_4 (.A0(rModDataWrite_15__N_1620[2]), .B0(rModDataWrite_15__N_1637[2]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[3]), 
          .B1(rModDataWrite_15__N_1637[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n14097), .COUT(n14098));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_4.INIT0 = 16'h5666;
    defparam add_320_4.INIT1 = 16'h5666;
    defparam add_320_4.INJECT1_0 = "NO";
    defparam add_320_4.INJECT1_1 = "NO";
    LUT4 i6873_2_lut (.A(PIC_DATA_IN_out_7), .B(PIC_WE_IN_c), .Z(data[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6873_2_lut.init = 16'h2222;
    CCU2D add_320_2 (.A0(rModDataWrite_15__N_1620[0]), .B0(rModDataWrite_15__N_1637[0]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1620[1]), 
          .B1(rModDataWrite_15__N_1637[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n14097));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_320_2.INIT0 = 16'h7000;
    defparam add_320_2.INIT1 = 16'h5666;
    defparam add_320_2.INJECT1_0 = "NO";
    defparam add_320_2.INJECT1_1 = "NO";
    CCU2D add_10506_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14289), 
          .S0(n2780));
    defparam add_10506_cout.INIT0 = 16'h0000;
    defparam add_10506_cout.INIT1 = 16'h0000;
    defparam add_10506_cout.INJECT1_0 = "NO";
    defparam add_10506_cout.INJECT1_1 = "NO";
    CCU2D add_10506_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14288), .COUT(n14289));
    defparam add_10506_21.INIT0 = 16'heeee;
    defparam add_10506_21.INIT1 = 16'heeee;
    defparam add_10506_21.INJECT1_0 = "NO";
    defparam add_10506_21.INJECT1_1 = "NO";
    CCU2D add_10506_19 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[17] ), .D0(n18264), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), .D1(lastAddress_31__N_1310), 
          .CIN(n14287), .COUT(n14288));
    defparam add_10506_19.INIT0 = 16'h00ce;
    defparam add_10506_19.INIT1 = 16'hff20;
    defparam add_10506_19.INJECT1_0 = "NO";
    defparam add_10506_19.INJECT1_1 = "NO";
    CCU2D add_10506_17 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n18271), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16] ), .D1(n18277), 
          .CIN(n14286), .COUT(n14287));
    defparam add_10506_17.INIT0 = 16'h00ce;
    defparam add_10506_17.INIT1 = 16'h00ce;
    defparam add_10506_17.INJECT1_0 = "NO";
    defparam add_10506_17.INJECT1_1 = "NO";
    CCU2D add_10506_15 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n18266), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n18262), 
          .CIN(n14285), .COUT(n14286));
    defparam add_10506_15.INIT0 = 16'h00ce;
    defparam add_10506_15.INIT1 = 16'h00ce;
    defparam add_10506_15.INJECT1_0 = "NO";
    defparam add_10506_15.INJECT1_1 = "NO";
    CCU2D add_10506_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n18273), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n18272), 
          .CIN(n14284), .COUT(n14285));
    defparam add_10506_13.INIT0 = 16'h00ce;
    defparam add_10506_13.INIT1 = 16'h00ce;
    defparam add_10506_13.INJECT1_0 = "NO";
    defparam add_10506_13.INJECT1_1 = "NO";
    CCU2D add_10506_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[9] ), .D0(n18268), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n18269), 
          .CIN(n14283), .COUT(n14284));
    defparam add_10506_11.INIT0 = 16'h00ce;
    defparam add_10506_11.INIT1 = 16'hff31;
    defparam add_10506_11.INJECT1_0 = "NO";
    defparam add_10506_11.INJECT1_1 = "NO";
    CCU2D add_10506_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[7] ), .D0(n18274), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), .D1(n18267), 
          .CIN(n14282), .COUT(n14283));
    defparam add_10506_9.INIT0 = 16'h00ce;
    defparam add_10506_9.INIT1 = 16'hff31;
    defparam add_10506_9.INJECT1_0 = "NO";
    defparam add_10506_9.INJECT1_1 = "NO";
    CCU2D add_10506_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[5] ), .D0(n18265), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[6] ), .D1(n18276), 
          .CIN(n14281), .COUT(n14282));
    defparam add_10506_7.INIT0 = 16'h00ce;
    defparam add_10506_7.INIT1 = 16'h00ce;
    defparam add_10506_7.INJECT1_0 = "NO";
    defparam add_10506_7.INJECT1_1 = "NO";
    CCU2D add_10506_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[3] ), .D0(n17409), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[4] ), .D1(n18275), 
          .CIN(n14280), .COUT(n14281));
    defparam add_10506_5.INIT0 = 16'h00ce;
    defparam add_10506_5.INIT1 = 16'h00ce;
    defparam add_10506_5.INJECT1_0 = "NO";
    defparam add_10506_5.INJECT1_1 = "NO";
    CCU2D add_10506_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[1] ), .D0(n17423), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[2] ), .D1(n18263), 
          .CIN(n14279), .COUT(n14280));
    defparam add_10506_3.INIT0 = 16'h00ce;
    defparam add_10506_3.INIT1 = 16'h00ce;
    defparam add_10506_3.INJECT1_0 = "NO";
    defparam add_10506_3.INJECT1_1 = "NO";
    CCU2D add_10506_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[0] ), 
          .D1(n18261), .COUT(n14279));
    defparam add_10506_1.INIT0 = 16'hF000;
    defparam add_10506_1.INIT1 = 16'h00ce;
    defparam add_10506_1.INJECT1_0 = "NO";
    defparam add_10506_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_265 (.A(n17444), .B(n17292), .C(n6105), .D(n17364), 
         .Z(LOGIC_CLOCK_enable_259)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    defparam i2_3_lut_4_lut_adj_265.init = 16'h0040;
    LUT4 i1_2_lut_adj_266 (.A(state_c[0]), .B(state[1]), .Z(n6105)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_adj_266.init = 16'h2222;
    LUT4 i1_4_lut_adj_267 (.A(n15454), .B(n17350), .C(state_c[5]), .D(n17445), 
         .Z(LOGIC_CLOCK_enable_251)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_267.init = 16'hccec;
    CCU2D lastAddress_18__I_0_0 (.A0(PIC_ADDR_IN_c_18), .B0(lastAddress[18]), 
          .C0(GND_net), .D0(GND_net), .A1(PIC_ADDR_IN_c_17), .B1(lastAddress[17]), 
          .C1(PIC_ADDR_IN_c_16), .D1(lastAddress[16]), .COUT(n13663));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[57:82])
    defparam lastAddress_18__I_0_0.INIT0 = 16'h9000;
    defparam lastAddress_18__I_0_0.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_0.INJECT1_0 = "NO";
    defparam lastAddress_18__I_0_0.INJECT1_1 = "YES";
    LUT4 i2_3_lut_adj_268 (.A(n15469), .B(state[4]), .C(state_c[3]), .Z(n15454)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut_adj_268.init = 16'h0808;
    CCU2D lastAddress_18__I_0_19 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n13667), .S0(BUS_DIRECTION_INTERNAL_N_1550));
    defparam lastAddress_18__I_0_19.INIT0 = 16'hFFFF;
    defparam lastAddress_18__I_0_19.INIT1 = 16'h0000;
    defparam lastAddress_18__I_0_19.INJECT1_0 = "NO";
    defparam lastAddress_18__I_0_19.INJECT1_1 = "NO";
    CCU2D lastAddress_18__I_0_19_10505 (.A0(PIC_ADDR_IN_c_3), .B0(lastAddress[3]), 
          .C0(PIC_ADDR_IN_c_2), .D0(lastAddress[2]), .A1(PIC_ADDR_IN_c_1), 
          .B1(lastAddress[1]), .C1(PIC_ADDR_IN_c_0), .D1(lastAddress[0]), 
          .CIN(n13666), .COUT(n13667));
    defparam lastAddress_18__I_0_19_10505.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_19_10505.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_19_10505.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_19_10505.INJECT1_1 = "YES";
    LUT4 i1_4_lut_adj_269 (.A(n15454), .B(n17350), .C(state_c[6]), .D(n15599), 
         .Z(LOGIC_CLOCK_enable_252)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_269.init = 16'hccec;
    LUT4 n16943_bdd_2_lut_4_lut (.A(state[1]), .B(n17389), .C(state_c[0]), 
         .D(n16943), .Z(state_7__N_1600[4])) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam n16943_bdd_2_lut_4_lut.init = 16'hff02;
    LUT4 i1_2_lut_4_lut (.A(state[1]), .B(n17389), .C(state_c[0]), .D(state_c[7]), 
         .Z(state_7__N_1600[7])) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_4_lut.init = 16'hff02;
    CCU2D lastAddress_18__I_0_17 (.A0(PIC_ADDR_IN_c_7), .B0(lastAddress[7]), 
          .C0(PIC_ADDR_IN_c_6), .D0(lastAddress[6]), .A1(PIC_ADDR_IN_c_5), 
          .B1(lastAddress[5]), .C1(PIC_ADDR_IN_c_4), .D1(lastAddress[4]), 
          .CIN(n13665), .COUT(n13666));
    defparam lastAddress_18__I_0_17.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_17.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_17.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_17.INJECT1_1 = "YES";
    LUT4 i2_3_lut_4_lut_adj_270 (.A(state[4]), .B(n17401), .C(n6105), 
         .D(state_c[3]), .Z(n15460)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i2_3_lut_4_lut_adj_270.init = 16'h0020;
    LUT4 i13045_3_lut_4_lut_4_lut (.A(n18260), .B(n63), .C(n2780), .D(BUS_VALID_N_1668), 
         .Z(LOGIC_CLOCK_enable_216)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i13045_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i11944_2_lut (.A(state_c[5]), .B(state_c[7]), .Z(n15599)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11944_2_lut.init = 16'heeee;
    LUT4 mux_725_i2_4_lut (.A(rModDataWrite[9]), .B(PIC_DATA_IN_out_1), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i2_4_lut.init = 16'h0aca;
    LUT4 mux_725_i3_4_lut (.A(rModDataWrite[10]), .B(PIC_DATA_IN_out_2), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i3_4_lut.init = 16'h0aca;
    LUT4 mux_725_i4_4_lut (.A(rModDataWrite[11]), .B(PIC_DATA_IN_out_3), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i4_4_lut.init = 16'h0aca;
    LUT4 mux_725_i5_4_lut (.A(rModDataWrite[12]), .B(PIC_DATA_IN_out_4), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i5_4_lut.init = 16'h0aca;
    LUT4 mux_725_i6_4_lut (.A(rModDataWrite[13]), .B(PIC_DATA_IN_out_5), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i6_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut (.A(n9), .B(\BUS_currGrantID[1] ), .C(n15657), .D(n17275), 
         .Z(LOGIC_CLOCK_enable_241)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i5_4_lut.init = 16'h0008;
    LUT4 mux_725_i7_4_lut (.A(rModDataWrite[14]), .B(PIC_DATA_IN_out_6), 
         .C(n15), .D(n5868), .Z(writeData_15__N_1719[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_725_i7_4_lut.init = 16'h0aca;
    LUT4 i6875_2_lut (.A(PIC_DATA_IN_out_9), .B(PIC_WE_IN_c), .Z(data[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6875_2_lut.init = 16'h2222;
    LUT4 i6876_2_lut (.A(PIC_DATA_IN_out_10), .B(PIC_WE_IN_c), .Z(data[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6876_2_lut.init = 16'h2222;
    LUT4 i11998_2_lut (.A(state_c[2]), .B(\BUS_currGrantID[0] ), .Z(n15657)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11998_2_lut.init = 16'heeee;
    LUT4 i6877_2_lut (.A(PIC_DATA_IN_out_11), .B(PIC_WE_IN_c), .Z(data[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6877_2_lut.init = 16'h2222;
    LUT4 i6878_2_lut (.A(PIC_DATA_IN_out_12), .B(PIC_WE_IN_c), .Z(data[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6878_2_lut.init = 16'h2222;
    LUT4 i6879_2_lut (.A(PIC_DATA_IN_out_13), .B(PIC_WE_IN_c), .Z(data[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6879_2_lut.init = 16'h2222;
    LUT4 i6880_2_lut (.A(PIC_DATA_IN_out_14), .B(PIC_WE_IN_c), .Z(data[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6880_2_lut.init = 16'h2222;
    LUT4 i6881_2_lut (.A(PIC_DATA_IN_out_15), .B(PIC_WE_IN_c), .Z(data[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i6881_2_lut.init = 16'h2222;
    LUT4 i13071_4_lut (.A(n17324), .B(n17292), .C(n15495), .D(n15), 
         .Z(LOGIC_CLOCK_enable_248)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;
    defparam i13071_4_lut.init = 16'h40c0;
    LUT4 i3_4_lut_adj_271 (.A(state[1]), .B(n15490), .C(state_c[3]), .D(n17364), 
         .Z(n15495)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_271.init = 16'hfffe;
    LUT4 i3850_3_lut (.A(LOGIC_CLOCK_enable_248), .B(n15), .C(n5868), 
         .Z(n7202)) /* synthesis lut_function=(A ((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i3850_3_lut.init = 16'ha2a2;
    LUT4 i1_2_lut_adj_272 (.A(state_c[0]), .B(state_c[2]), .Z(n15490)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_272.init = 16'heeee;
    CCU2D add_10511_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n14177), 
          .S0(BUS_VALID_N_1668));
    defparam add_10511_cout.INIT0 = 16'h0000;
    defparam add_10511_cout.INIT1 = 16'h0000;
    defparam add_10511_cout.INJECT1_0 = "NO";
    defparam add_10511_cout.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_273 (.A(state_c[0]), .B(n17444), .C(state[1]), .D(n17363), 
         .Z(n15)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i3_4_lut_adj_273.init = 16'hffef;
    CCU2D add_10511_13 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n14176), .COUT(n14177));
    defparam add_10511_13.INIT0 = 16'heeee;
    defparam add_10511_13.INIT1 = 16'heeee;
    defparam add_10511_13.INJECT1_0 = "NO";
    defparam add_10511_13.INJECT1_1 = "NO";
    LUT4 readData_15__I_0_i2_4_lut (.A(transferMode[1]), .B(writeData_c[1]), 
         .C(n9950), .D(n63), .Z(\BUS_DATA_INTERNAL[1] )) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(68[23:106])
    defparam readData_15__I_0_i2_4_lut.init = 16'h0cac;
    LUT4 readData_15__I_0_i3_4_lut (.A(transferMode[2]), .B(writeData_c[2]), 
         .C(n9950), .D(n63), .Z(\BUS_DATA_INTERNAL[2] )) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(68[23:106])
    defparam readData_15__I_0_i3_4_lut.init = 16'h0cac;
    CCU2D add_10511_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[17] ), .D0(n18264), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), .D1(lastAddress_31__N_1310), 
          .CIN(n14175), .COUT(n14176));
    defparam add_10511_11.INIT0 = 16'h00ce;
    defparam add_10511_11.INIT1 = 16'hff20;
    defparam add_10511_11.INJECT1_0 = "NO";
    defparam add_10511_11.INJECT1_1 = "NO";
    PFUMX i13410 (.BLUT(n17474), .ALUT(n17475), .C0(state_c[0]), .Z(state_7__N_1600[0]));
    LUT4 readData_15__I_0_i4_4_lut (.A(transferMode[3]), .B(writeData_c[3]), 
         .C(n9950), .D(n63), .Z(\BUS_DATA_INTERNAL[3] )) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(68[23:106])
    defparam readData_15__I_0_i4_4_lut.init = 16'h0cac;
    CCU2D add_10511_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n18271), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16] ), .D1(n18277), 
          .CIN(n14174), .COUT(n14175));
    defparam add_10511_9.INIT0 = 16'h00ce;
    defparam add_10511_9.INIT1 = 16'h00ce;
    defparam add_10511_9.INJECT1_0 = "NO";
    defparam add_10511_9.INJECT1_1 = "NO";
    LUT4 n6241_bdd_3_lut_13373_4_lut (.A(n17444), .B(n17401), .C(state[4]), 
         .D(state_c[0]), .Z(n16941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    defparam n6241_bdd_3_lut_13373_4_lut.init = 16'hf0e0;
    LUT4 i2_3_lut_rep_342_4_lut (.A(n17444), .B(n17401), .C(state_c[0]), 
         .D(state[1]), .Z(n17350)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    defparam i2_3_lut_rep_342_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_4_lut_adj_274 (.A(state_c[5]), .B(n17445), .C(state_c[3]), 
         .D(n15490), .Z(n15491)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_274.init = 16'hfffe;
    CCU2D add_10511_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n18266), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n18262), 
          .CIN(n14173), .COUT(n14174));
    defparam add_10511_7.INIT0 = 16'h00ce;
    defparam add_10511_7.INIT1 = 16'h00ce;
    defparam add_10511_7.INJECT1_0 = "NO";
    defparam add_10511_7.INJECT1_1 = "NO";
    CCU2D lastAddress_18__I_0_15 (.A0(PIC_ADDR_IN_c_11), .B0(lastAddress[11]), 
          .C0(PIC_ADDR_IN_c_10), .D0(lastAddress[10]), .A1(PIC_ADDR_IN_c_9), 
          .B1(lastAddress[9]), .C1(PIC_ADDR_IN_c_8), .D1(lastAddress[8]), 
          .CIN(n13664), .COUT(n13665));
    defparam lastAddress_18__I_0_15.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_15.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_15.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_15.INJECT1_1 = "YES";
    CCU2D lastAddress_18__I_0_13 (.A0(PIC_ADDR_IN_c_15), .B0(lastAddress[15]), 
          .C0(PIC_ADDR_IN_c_14), .D0(lastAddress[14]), .A1(PIC_ADDR_IN_c_13), 
          .B1(lastAddress[13]), .C1(PIC_ADDR_IN_c_12), .D1(lastAddress[12]), 
          .CIN(n13663), .COUT(n13664));
    defparam lastAddress_18__I_0_13.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_13.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_13.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_13.INJECT1_1 = "YES";
    LUT4 i11923_2_lut_3_lut_4_lut (.A(state[1]), .B(n17444), .C(n17401), 
         .D(state[4]), .Z(n15577)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i11923_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_316_3_lut_4_lut (.A(state[1]), .B(n17444), .C(n17401), 
         .D(state[4]), .Z(n17324)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_316_3_lut_4_lut.init = 16'hfffe;
    PFUMX i13231 (.BLUT(n16942), .ALUT(n16941), .C0(state[1]), .Z(n16943));
    LUT4 i1_4_lut_adj_275 (.A(n17350), .B(state_c[0]), .C(n12), .D(n15577), 
         .Z(BUS_REQ_N_1761)) /* synthesis lut_function=(A+(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_275.init = 16'hfafb;
    LUT4 i1_4_lut_adj_276 (.A(\BUS_req[2] ), .B(state[4]), .C(n6_adj_1879), 
         .D(n17389), .Z(n12)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_276.init = 16'haaa2;
    LUT4 i2_4_lut_adj_277 (.A(state[1]), .B(n17390), .C(n17434), .D(n17270), 
         .Z(n6_adj_1879)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;
    defparam i2_4_lut_adj_277.init = 16'haaba;
    
endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 00:39:41 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 76 -num_rows 512 -rdata_width 76 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr76951276951211d16619 -pmi -lang verilog  */
/* Tue Jan 12 00:39:40 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr76951276951211d16619 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [75:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [75:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(scuba_vlo), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(), .DO12(Q[75]), 
        .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), .DO8(), .DO7(), .DO6(), 
        .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_0_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_1_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_2_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_3_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr76951276951211d16619__PMIP__512__76__76B
    // exemplar attribute pmi_ram_dpXbnonesadr76951276951211d16619_0_4_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 00:42:54 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 113 -num_rows 512 -rdata_width 113 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1139512113951211f50d4a -pmi -lang verilog  */
/* Tue Jan 12 00:42:53 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1139512113951211f50d4a (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [112:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [112:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(Q[112]), 
        .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), .DO8(), 
        .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 00:51:26 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 113 -num_rows 512 -rdata_width 113 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1139512113951211f50d4a -pmi -lang verilog  */
/* Tue Jan 12 00:51:25 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1139512113951211f50d4a (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [112:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [112:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(Q[112]), 
        .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), .DO8(), 
        .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 00:54:49 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 129 -num_rows 512 -rdata_width 129 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1299512129951211f54899 -pmi -lang verilog  */
/* Tue Jan 12 00:54:48 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1299512129951211f54899 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [128:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [128:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(scuba_vlo), .DI3(scuba_vlo), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(), .DO12(), 
        .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), .DO8(), .DO7(), .DO6(), 
        .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_0_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_1_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_2_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_3_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_4_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_5_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_6_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1299512129951211f54899__PMIP__512__129__129B
    // exemplar attribute pmi_ram_dpXbnonesadr1299512129951211f54899_0_7_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:00:09 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 175 -num_rows 512 -rdata_width 175 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1759512175951211f54f9f -pmi -lang verilog  */
/* Tue Jan 12 01:00:08 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1759512175951211f54f9f (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [174:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [174:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(Data[174]), .DI11(Data[173]), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(Q[174]), .DO2(Q[173]), 
        .DO1(Q[172]), .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:07:33 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 175 -num_rows 512 -rdata_width 175 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1759512175951211f54f9f -pmi -lang verilog  */
/* Tue Jan 12 01:07:32 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1759512175951211f54f9f (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [174:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [174:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(Data[174]), .DI11(Data[173]), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(Q[174]), .DO2(Q[173]), 
        .DO1(Q[172]), .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:13:18 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 175 -num_rows 512 -rdata_width 175 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1759512175951211f54f9f -pmi -lang verilog  */
/* Tue Jan 12 01:13:17 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1759512175951211f54f9f (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [174:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [174:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(Data[174]), .DI11(Data[173]), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(Q[174]), .DO2(Q[173]), 
        .DO1(Q[172]), .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:22:40 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 175 -num_rows 512 -rdata_width 175 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1759512175951211f54f9f -pmi -lang verilog  */
/* Tue Jan 12 01:22:39 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1759512175951211f54f9f (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [174:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [174:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(Data[174]), .DI11(Data[173]), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(Q[174]), .DO2(Q[173]), 
        .DO1(Q[172]), .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:26:48 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 175 -num_rows 512 -rdata_width 175 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1759512175951211f54f9f -pmi -lang verilog  */
/* Tue Jan 12 01:26:47 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1759512175951211f54f9f (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [174:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [174:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(Data[174]), .DI11(Data[173]), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(Q[174]), .DO2(Q[173]), 
        .DO1(Q[172]), .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:30:01 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 175 -num_rows 512 -rdata_width 175 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1759512175951211f54f9f -pmi -lang verilog  */
/* Tue Jan 12 01:30:00 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1759512175951211f54f9f (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [174:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [174:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(Data[174]), .DI11(Data[173]), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(Q[174]), .DO2(Q[173]), 
        .DO1(Q[172]), .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1759512175951211f54f9f__PMIP__512__175__175B
    // exemplar attribute pmi_ram_dpXbnonesadr1759512175951211f54f9f_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:34:01 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 113 -num_rows 512 -rdata_width 113 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1139512113951211f50d4a -pmi -lang verilog  */
/* Tue Jan 12 01:34:00 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1139512113951211f50d4a (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [112:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [112:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(Q[112]), 
        .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), .DO8(), 
        .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_0_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_1_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_2_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_3_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_4_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_5_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1139512113951211f50d4a__PMIP__512__113__113B
    // exemplar attribute pmi_ram_dpXbnonesadr1139512113951211f50d4a_0_6_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:36:49 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 148 -num_rows 512 -rdata_width 148 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1489512148951211f54e2b -pmi -lang verilog  */
/* Tue Jan 12 01:36:48 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1489512148951211f54e2b (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [147:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [147:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(scuba_vlo), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(), .DO12(Q[147]), 
        .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), .DO8(), .DO7(), .DO6(), 
        .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_0_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_1_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_2_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_3_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_4_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_5_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_6_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_7_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1489512148951211f54e2b__PMIP__512__148__148B
    // exemplar attribute pmi_ram_dpXbnonesadr1489512148951211f54e2b_0_8_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:40:27 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 111 -num_rows 512 -rdata_width 111 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1119512111951211f4fc04 -pmi -lang verilog  */
/* Tue Jan 12 01:40:26 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1119512111951211f4fc04 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [110:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [110:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(scuba_vlo), .DI9(scuba_vlo), 
        .DI8(scuba_vlo), .DI7(scuba_vlo), .DI6(scuba_vlo), .DI5(scuba_vlo), 
        .DI4(scuba_vlo), .DI3(scuba_vlo), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(), .DO16(), .DO15(), .DO14(), .DO13(), .DO12(), 
        .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), .DO8(), .DO7(), .DO6(), 
        .DO5(), .DO4(), .DO3(), .DO2(), .DO1(), .DO0())
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_0_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_1_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_2_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_3_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_4_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_5_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1119512111951211f4fc04__PMIP__512__111__111B
    // exemplar attribute pmi_ram_dpXbnonesadr1119512111951211f4fc04_0_6_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 01:45:01 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 143 -num_rows 512 -rdata_width 143 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1439512143951211f525f7 -pmi -lang verilog  */
/* Tue Jan 12 01:45:00 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1439512143951211f525f7 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [142:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [142:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0 (.DI17(scuba_vlo), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_0_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_1_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_2_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_3_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_4_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_5_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_6_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1439512143951211f525f7__PMIP__512__143__143B
    // exemplar attribute pmi_ram_dpXbnonesadr1439512143951211f525f7_0_7_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 11:55:15 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 11:55:14 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 12:01:09 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 12:01:08 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 12:04:51 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 12:04:50 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 12:09:44 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 12:09:44 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 12:12:34 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 12:12:33 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 12:20:42 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 12:20:41 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 16 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner24168de3ddc -pmi -lang verilog  */
/* Tue Jan 12 12:24:11 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner24168de3ddc (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [3:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [3:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire dataout1_ffin;
    wire dataout0_ffin;
    wire dec0_wre3;
    wire scuba_vhi;

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(scuba_vhi), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(dataout0_ffin), .DO1(dataout1_ffin), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B" */
             /* synthesis COMP="mem_0_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner24168de3ddc__PMI__16__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 173 -num_rows 512 -rdata_width 173 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr1739512173951211f540e2 -pmi -lang verilog  */
/* Tue Jan 12 12:24:10 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr1739512173951211f540e2 (WrAddress, RdAddress, 
    Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [8:0] WrAddress;
    input wire [8:0] RdAddress;
    input wire [172:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [172:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 (.DI17(Data[17]), 
        .DI16(Data[16]), .DI15(Data[15]), .DI14(Data[14]), .DI13(Data[13]), 
        .DI12(Data[12]), .DI11(Data[11]), .DI10(Data[10]), .DI9(Data[9]), 
        .DI8(Data[8]), .DI7(Data[7]), .DI6(Data[6]), .DI5(Data[5]), .DI4(Data[4]), 
        .DI3(Data[3]), .DI2(Data[2]), .DI1(Data[1]), .DI0(Data[0]), .ADW8(WrAddress[8]), 
        .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), 
        .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), 
        .BE1(scuba_vhi), .BE0(scuba_vhi), .CEW(WrClockEn), .CLKW(WrClock), 
        .CSW2(scuba_vlo), .CSW1(scuba_vlo), .CSW0(WE), .ADR12(RdAddress[8]), 
        .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), .ADR9(RdAddress[5]), 
        .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), .ADR5(RdAddress[1]), 
        .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), .ADR1(scuba_vlo), 
        .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), .CLKR(RdClock), 
        .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), .RST(Reset), 
        .DO17(Q[8]), .DO16(Q[7]), .DO15(Q[6]), .DO14(Q[5]), .DO13(Q[4]), 
        .DO12(Q[3]), .DO11(Q[2]), .DO10(Q[1]), .DO9(Q[0]), .DO8(Q[17]), 
        .DO7(Q[16]), .DO6(Q[15]), .DO5(Q[14]), .DO4(Q[13]), .DO3(Q[12]), 
        .DO2(Q[11]), .DO1(Q[10]), .DO0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 (.DI17(Data[35]), 
        .DI16(Data[34]), .DI15(Data[33]), .DI14(Data[32]), .DI13(Data[31]), 
        .DI12(Data[30]), .DI11(Data[29]), .DI10(Data[28]), .DI9(Data[27]), 
        .DI8(Data[26]), .DI7(Data[25]), .DI6(Data[24]), .DI5(Data[23]), 
        .DI4(Data[22]), .DI3(Data[21]), .DI2(Data[20]), .DI1(Data[19]), 
        .DI0(Data[18]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[26]), .DO16(Q[25]), .DO15(Q[24]), .DO14(Q[23]), 
        .DO13(Q[22]), .DO12(Q[21]), .DO11(Q[20]), .DO10(Q[19]), .DO9(Q[18]), 
        .DO8(Q[35]), .DO7(Q[34]), .DO6(Q[33]), .DO5(Q[32]), .DO4(Q[31]), 
        .DO3(Q[30]), .DO2(Q[29]), .DO1(Q[28]), .DO0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 (.DI17(Data[53]), 
        .DI16(Data[52]), .DI15(Data[51]), .DI14(Data[50]), .DI13(Data[49]), 
        .DI12(Data[48]), .DI11(Data[47]), .DI10(Data[46]), .DI9(Data[45]), 
        .DI8(Data[44]), .DI7(Data[43]), .DI6(Data[42]), .DI5(Data[41]), 
        .DI4(Data[40]), .DI3(Data[39]), .DI2(Data[38]), .DI1(Data[37]), 
        .DI0(Data[36]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[44]), .DO16(Q[43]), .DO15(Q[42]), .DO14(Q[41]), 
        .DO13(Q[40]), .DO12(Q[39]), .DO11(Q[38]), .DO10(Q[37]), .DO9(Q[36]), 
        .DO8(Q[53]), .DO7(Q[52]), .DO6(Q[51]), .DO5(Q[50]), .DO4(Q[49]), 
        .DO3(Q[48]), .DO2(Q[47]), .DO1(Q[46]), .DO0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 (.DI17(Data[71]), 
        .DI16(Data[70]), .DI15(Data[69]), .DI14(Data[68]), .DI13(Data[67]), 
        .DI12(Data[66]), .DI11(Data[65]), .DI10(Data[64]), .DI9(Data[63]), 
        .DI8(Data[62]), .DI7(Data[61]), .DI6(Data[60]), .DI5(Data[59]), 
        .DI4(Data[58]), .DI3(Data[57]), .DI2(Data[56]), .DI1(Data[55]), 
        .DI0(Data[54]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[62]), .DO16(Q[61]), .DO15(Q[60]), .DO14(Q[59]), 
        .DO13(Q[58]), .DO12(Q[57]), .DO11(Q[56]), .DO10(Q[55]), .DO9(Q[54]), 
        .DO8(Q[71]), .DO7(Q[70]), .DO6(Q[69]), .DO5(Q[68]), .DO4(Q[67]), 
        .DO3(Q[66]), .DO2(Q[65]), .DO1(Q[64]), .DO0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 (.DI17(Data[89]), 
        .DI16(Data[88]), .DI15(Data[87]), .DI14(Data[86]), .DI13(Data[85]), 
        .DI12(Data[84]), .DI11(Data[83]), .DI10(Data[82]), .DI9(Data[81]), 
        .DI8(Data[80]), .DI7(Data[79]), .DI6(Data[78]), .DI5(Data[77]), 
        .DI4(Data[76]), .DI3(Data[75]), .DI2(Data[74]), .DI1(Data[73]), 
        .DI0(Data[72]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[80]), .DO16(Q[79]), .DO15(Q[78]), .DO14(Q[77]), 
        .DO13(Q[76]), .DO12(Q[75]), .DO11(Q[74]), .DO10(Q[73]), .DO9(Q[72]), 
        .DO8(Q[89]), .DO7(Q[88]), .DO6(Q[87]), .DO5(Q[86]), .DO4(Q[85]), 
        .DO3(Q[84]), .DO2(Q[83]), .DO1(Q[82]), .DO0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 (.DI17(Data[107]), 
        .DI16(Data[106]), .DI15(Data[105]), .DI14(Data[104]), .DI13(Data[103]), 
        .DI12(Data[102]), .DI11(Data[101]), .DI10(Data[100]), .DI9(Data[99]), 
        .DI8(Data[98]), .DI7(Data[97]), .DI6(Data[96]), .DI5(Data[95]), 
        .DI4(Data[94]), .DI3(Data[93]), .DI2(Data[92]), .DI1(Data[91]), 
        .DI0(Data[90]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[98]), .DO16(Q[97]), .DO15(Q[96]), .DO14(Q[95]), 
        .DO13(Q[94]), .DO12(Q[93]), .DO11(Q[92]), .DO10(Q[91]), .DO9(Q[90]), 
        .DO8(Q[107]), .DO7(Q[106]), .DO6(Q[105]), .DO5(Q[104]), .DO4(Q[103]), 
        .DO3(Q[102]), .DO2(Q[101]), .DO1(Q[100]), .DO0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 (.DI17(Data[125]), 
        .DI16(Data[124]), .DI15(Data[123]), .DI14(Data[122]), .DI13(Data[121]), 
        .DI12(Data[120]), .DI11(Data[119]), .DI10(Data[118]), .DI9(Data[117]), 
        .DI8(Data[116]), .DI7(Data[115]), .DI6(Data[114]), .DI5(Data[113]), 
        .DI4(Data[112]), .DI3(Data[111]), .DI2(Data[110]), .DI1(Data[109]), 
        .DI0(Data[108]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[116]), .DO16(Q[115]), .DO15(Q[114]), .DO14(Q[113]), 
        .DO13(Q[112]), .DO12(Q[111]), .DO11(Q[110]), .DO10(Q[109]), .DO9(Q[108]), 
        .DO8(Q[125]), .DO7(Q[124]), .DO6(Q[123]), .DO5(Q[122]), .DO4(Q[121]), 
        .DO3(Q[120]), .DO2(Q[119]), .DO1(Q[118]), .DO0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 (.DI17(Data[143]), 
        .DI16(Data[142]), .DI15(Data[141]), .DI14(Data[140]), .DI13(Data[139]), 
        .DI12(Data[138]), .DI11(Data[137]), .DI10(Data[136]), .DI9(Data[135]), 
        .DI8(Data[134]), .DI7(Data[133]), .DI6(Data[132]), .DI5(Data[131]), 
        .DI4(Data[130]), .DI3(Data[129]), .DI2(Data[128]), .DI1(Data[127]), 
        .DI0(Data[126]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[134]), .DO16(Q[133]), .DO15(Q[132]), .DO14(Q[131]), 
        .DO13(Q[130]), .DO12(Q[129]), .DO11(Q[128]), .DO10(Q[127]), .DO9(Q[126]), 
        .DO8(Q[143]), .DO7(Q[142]), .DO6(Q[141]), .DO5(Q[140]), .DO4(Q[139]), 
        .DO3(Q[138]), .DO2(Q[137]), .DO1(Q[136]), .DO0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 (.DI17(Data[161]), 
        .DI16(Data[160]), .DI15(Data[159]), .DI14(Data[158]), .DI13(Data[157]), 
        .DI12(Data[156]), .DI11(Data[155]), .DI10(Data[154]), .DI9(Data[153]), 
        .DI8(Data[152]), .DI7(Data[151]), .DI6(Data[150]), .DI5(Data[149]), 
        .DI4(Data[148]), .DI3(Data[147]), .DI2(Data[146]), .DI1(Data[145]), 
        .DI0(Data[144]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[152]), .DO16(Q[151]), .DO15(Q[150]), .DO14(Q[149]), 
        .DO13(Q[148]), .DO12(Q[147]), .DO11(Q[146]), .DO10(Q[145]), .DO9(Q[144]), 
        .DO8(Q[161]), .DO7(Q[160]), .DO6(Q[159]), .DO5(Q[158]), .DO4(Q[157]), 
        .DO3(Q[156]), .DO2(Q[155]), .DO1(Q[154]), .DO0(Q[153]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_R = "0b000" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.CSDECODE_W = "0b001" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.REGMODE = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_R = 18 ;
    defparam pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0.DATA_WIDTH_W = 18 ;
    PDPW8KC pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 (.DI17(scuba_vlo), 
        .DI16(scuba_vlo), .DI15(scuba_vlo), .DI14(scuba_vlo), .DI13(scuba_vlo), 
        .DI12(scuba_vlo), .DI11(scuba_vlo), .DI10(Data[172]), .DI9(Data[171]), 
        .DI8(Data[170]), .DI7(Data[169]), .DI6(Data[168]), .DI5(Data[167]), 
        .DI4(Data[166]), .DI3(Data[165]), .DI2(Data[164]), .DI1(Data[163]), 
        .DI0(Data[162]), .ADW8(WrAddress[8]), .ADW7(WrAddress[7]), .ADW6(WrAddress[6]), 
        .ADW5(WrAddress[5]), .ADW4(WrAddress[4]), .ADW3(WrAddress[3]), .ADW2(WrAddress[2]), 
        .ADW1(WrAddress[1]), .ADW0(WrAddress[0]), .BE1(scuba_vhi), .BE0(scuba_vhi), 
        .CEW(WrClockEn), .CLKW(WrClock), .CSW2(scuba_vlo), .CSW1(scuba_vlo), 
        .CSW0(WE), .ADR12(RdAddress[8]), .ADR11(RdAddress[7]), .ADR10(RdAddress[6]), 
        .ADR9(RdAddress[5]), .ADR8(RdAddress[4]), .ADR7(RdAddress[3]), .ADR6(RdAddress[2]), 
        .ADR5(RdAddress[1]), .ADR4(RdAddress[0]), .ADR3(scuba_vlo), .ADR2(scuba_vlo), 
        .ADR1(scuba_vlo), .ADR0(scuba_vlo), .CER(RdClockEn), .OCER(RdClockEn), 
        .CLKR(RdClock), .CSR2(scuba_vlo), .CSR1(scuba_vlo), .CSR0(scuba_vlo), 
        .RST(Reset), .DO17(Q[170]), .DO16(Q[169]), .DO15(Q[168]), .DO14(Q[167]), 
        .DO13(Q[166]), .DO12(Q[165]), .DO11(Q[164]), .DO10(Q[163]), .DO9(Q[162]), 
        .DO8(), .DO7(), .DO6(), .DO5(), .DO4(), .DO3(), .DO2(), .DO1(Q[172]), 
        .DO0(Q[171]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_0_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_1_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_2_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_3_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_4_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_5_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_6_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_7_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_8_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr1739512173951211f540e2__PMIP__512__173__173B
    // exemplar attribute pmi_ram_dpXbnonesadr1739512173951211f540e2_0_9_0 MEM_INIT_FILE 
    // exemplar end

endmodule
