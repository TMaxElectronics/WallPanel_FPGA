// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Sun Jan 10 17:24:40 2021
//
// Verilog Description of module Master
//

module Master (CLK, UART_RX, UART_TX, Matrix_DATA_Out, Matrix_LINE_SEL_Out, 
            Matrix_CTRL_Out, SRAM_OE, SRAM_WE, SRAM_CE, SRAM_DATA, 
            SRAM_ADDR, PIC_OE, PIC_WE_IN, PIC_CS, PIC_ADDR_IN, PIC_DATA_IN, 
            PIC_READY, LED);   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(6[8:14])
    input CLK;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    input UART_RX;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(10[3:10])
    output UART_TX;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(11[3:10])
    output [11:0]Matrix_DATA_Out;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    output [3:0]Matrix_LINE_SEL_Out;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    output [2:0]Matrix_CTRL_Out;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    output SRAM_OE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(17[3:10])
    output SRAM_WE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(18[3:10])
    output SRAM_CE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(19[3:10])
    inout [15:0]SRAM_DATA;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(20[3:12])
    output [17:0]SRAM_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    input PIC_OE;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(23[3:9])
    input PIC_WE_IN;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    input PIC_CS;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(25[3:9])
    input [18:0]PIC_ADDR_IN;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    inout [15:0]PIC_DATA_IN;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(27[3:14])
    output PIC_READY;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(28[3:12])
    output [7:0]LED;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    
    wire CLK_c /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    wire PIXEL_CLOCK /* synthesis SET_AS_NETWORK=PIXEL_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(43[8:19])
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(90[8:15])
    wire PIXEL_CLOCK_N_302 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(82[9:22])
    wire LOGIC_CLOCK_N_116 /* synthesis is_clock=1, is_inv_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(73[9:17])
    
    wire GND_net, VCC_net, Matrix_DATA_Out_c_11, Matrix_DATA_Out_c_10, 
        Matrix_DATA_Out_c_9, Matrix_DATA_Out_c_8, Matrix_DATA_Out_c_7, 
        Matrix_DATA_Out_c_6, Matrix_DATA_Out_c_5, Matrix_DATA_Out_c_4, 
        Matrix_DATA_Out_c_3, Matrix_DATA_Out_c_2, Matrix_DATA_Out_c_1, 
        Matrix_DATA_Out_c_0, Matrix_LINE_SEL_Out_c_2, Matrix_LINE_SEL_Out_c_1, 
        Matrix_LINE_SEL_Out_c_0, Matrix_CTRL_Out_c_2, Matrix_CTRL_Out_c_1, 
        Matrix_CTRL_Out_c_0, SRAM_OE_c, SRAM_WE_c, n10855, SRAM_ADDR_c_17, 
        SRAM_ADDR_c_16, SRAM_ADDR_c_15, SRAM_ADDR_c_14, SRAM_ADDR_c_13, 
        SRAM_ADDR_c_12, SRAM_ADDR_c_11, SRAM_ADDR_c_10, SRAM_ADDR_c_9, 
        SRAM_ADDR_c_8, SRAM_ADDR_c_7, SRAM_ADDR_c_6, SRAM_ADDR_c_5, 
        SRAM_ADDR_c_4, SRAM_ADDR_c_3, SRAM_ADDR_c_2, SRAM_ADDR_c_1, 
        SRAM_ADDR_c_0, PIC_OE_c, PIC_WE_IN_c, PIC_ADDR_IN_c_18, PIC_ADDR_IN_c_17, 
        PIC_ADDR_IN_c_16, PIC_ADDR_IN_c_15, PIC_ADDR_IN_c_14, PIC_ADDR_IN_c_13, 
        PIC_ADDR_IN_c_12, PIC_ADDR_IN_c_11, PIC_ADDR_IN_c_10, PIC_ADDR_IN_c_9, 
        PIC_ADDR_IN_c_8, PIC_ADDR_IN_c_7, PIC_ADDR_IN_c_6, PIC_ADDR_IN_c_5, 
        PIC_ADDR_IN_c_4, PIC_ADDR_IN_c_3, PIC_ADDR_IN_c_2, PIC_ADDR_IN_c_1, 
        PIC_ADDR_IN_c_0, PIC_READY_c;
    wire [15:0]BUS_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(48[8:16])
    wire [31:0]BUS_addr;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    
    wire BUS_DONE;
    wire [3:0]BUS_req;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(54[8:15])
    wire [3:0]BUS_currGrantID;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    wire [15:0]PIC_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(58[8:16])
    
    wire n54, n37, n3244, n3245, n3246;
    wire [15:0]MATRIX_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(69[8:19])
    wire [15:0]MDM_data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(73[8:16])
    
    wire n3360, n3152, n3151, n3150, n3149, MDM_done, BUS_DONE_OVERRIDE;
    wire [7:0]VRAM_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(88[8:17])
    wire [9:0]n3028;
    wire [9:0]n3027;
    wire [9:0]VRAM_DATA;
    wire [9:0]n3031;
    wire [9:0]n3030;
    wire [9:0]n3029;
    wire [9:0]n3037;
    wire [9:0]n3036;
    wire [9:0]n3035;
    wire [9:0]n3034;
    wire [9:0]n3033;
    wire [9:0]n3032;
    wire [4:0]MATRIX_CURRROW;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(91[8:22])
    
    wire n34, n60, n42, n71, n7, BUS_currGrantID_3__N_54, n3234, 
        n3233, n3232, n3231, n3238, n3237, n3236, n3235, n3240, 
        n3239;
    wire [3:0]BUS_currGrantID_3__N_72;
    
    wire n11153, n11193;
    wire [15:0]\PWMArray[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(73[9:17])
    
    wire n5648, n33, n11152, n3354, n11151, n3359, n3358, n45, 
        n64, n62, n61, n59, n56, n46, n4545, n3169, n3168, 
        n3167, n3166, n3165, n3164, n3163, n3162, n3161, n3160, 
        n3159, n11331, n11206, n11222, n3353, n3355, n3365, n3364, 
        n11101, n11108, n3349, n3361, n3371, n5, n3375, n52, 
        n3363, LOGIC_CLOCK_enable_71, n87;
    wire [15:0]currPWMCount;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(86[9:21])
    wire [15:0]currPWMCountMax;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(87[9:24])
    
    wire n3170, n2025, WRITE_DONE, n3370, n3351, n58, n48, n1184, 
        n4537, n57, n3377, n3372, n43, n3314, n3380, n3374, 
        n3373, n3357, SRAM_DATA_out_13, n6, BUS_VALID_N_113, PWMArray_0__12__N_110;
    wire [4:0]currReadRow;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(54[9:20])
    wire [4:0]lastReadRow;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(55[9:20])
    wire [7:0]xOffset;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(62[9:16])
    wire [7:0]yOffset;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(63[9:16])
    wire [31:0]BUS_ADDR_INTERNAL;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(81[9:26])
    
    wire n11334;
    wire [15:0]otherData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(97[9:18])
    
    wire reset, n11333;
    wire [15:0]BUS_DATA_INTERNAL_adj_1354;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(104[9:26])
    wire [9:0]GR_WR_DOUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(133[9:19])
    wire [7:0]GR_WR_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(136[9:19])
    
    wire n10349, n3367, n2259, n2260, n2261, n2262, n2263, n2264, 
        n2265, n2266, n3315, n3316, n3317, n3318, n3319, n3320, 
        n3321, n3322, n3323, n3324, n11332, n3325, n3326, n3327, 
        n3328, n3329, n11146, n11004, n3330, n3272, n3273, n3274, 
        n11145, n3275, n3277, n3278, n11144, n11139, n11138, n11137, 
        n3379, n47, n49, n11327, n36, n11326, n3350, n11132, 
        n11131, n3356, n11130, n11325, n7167, n3331, n3332, n3333, 
        n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
        n3342, n3343, n3344, n41, n1921, n3144, n3143, n3142, 
        n3141, n3140, n3139, n39, n13158, n11012, n13157, n11125, 
        n11124, n11123, n3135, n3134, n3133, n3132, n3131, n3130, 
        n3129, n3128, n3127, n3126, n3125, n3124, n3123, n3122, 
        n3121, n13156, n3213, n3212, n3211, n3210, n3209, n13155, 
        BUS_DONE_OUT_N_626, n4, n3247, n3248, n3249, n13154, n12219, 
        n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, 
        n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, 
        n3266, n3267, n3268, n3269, n5_adj_1307, n3270, n3271, 
        n1886, n13153, n13152, n3366, n3345, n2589, n3104, n11118, 
        n3105, n3106, n3107, n3108, n13151, n4541, n55, n7_adj_1308, 
        n12218, n63, n10350, n2198;
    wire [31:0]lastAddress;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(29[8:19])
    wire [15:0]BUS_DATA_INTERNAL_adj_1362;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(30[8:25])
    
    wire BUS_DONE_INTERNAL, lastAddress_31__N_778, lastAddress_31__N_845, 
        lastAddress_31__N_863, lastAddress_31__N_783, lastAddress_31__N_860, 
        lastAddress_31__N_782, lastAddress_31__N_857, lastAddress_31__N_781, 
        lastAddress_31__N_854, lastAddress_31__N_780, lastAddress_31__N_851, 
        lastAddress_31__N_779, lastAddress_31__N_848, lastAddress_31__N_884, 
        lastAddress_31__N_790, SRAM_WE_N_704, n4_adj_1313, n4_adj_1314, 
        n13150, n13149, n13148, n40, n11117, n12348, n13147, n3352, 
        n12344, n12342, n13146, n13145, n13144, n3109, n3110, 
        n3111, n3112, n3113, n6_adj_1315, n11116, n13143, lastAddress_31__N_760, 
        lastAddress_31__N_777, lastAddress_31__N_842, lastAddress_31__N_776, 
        lastAddress_31__N_839, lastAddress_31__N_775, lastAddress_31__N_836, 
        lastAddress_31__N_774, lastAddress_31__N_833, lastAddress_31__N_773, 
        lastAddress_31__N_830, lastAddress_31__N_827, lastAddress_31__N_881, 
        lastAddress_31__N_789, lastAddress_31__N_878, lastAddress_31__N_788, 
        lastAddress_31__N_875, lastAddress_31__N_787, lastAddress_31__N_872, 
        lastAddress_31__N_786, lastAddress_31__N_869, lastAddress_31__N_785, 
        lastAddress_31__N_866, lastAddress_31__N_784, BUS_DIRECTION_INTERNAL;
    wire [15:0]BUS_DATA_INTERNAL_adj_1373;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(39[8:25])
    wire [31:0]BUS_ADDR_INTERNAL_adj_1374;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(40[8:25])
    
    wire WRITE_DONE_adj_1337;
    wire [15:0]writeData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(46[8:17])
    wire [7:0]state_adj_1377;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    
    wire BUS_VALID_N_1118, n12332, transferMode_3__N_1115, n3114, n3115, 
        n12217, n5045, n12329, n3153, n13142, n13141, n13140, 
        n3116, n13139;
    wire [7:0]state_7__N_1050;
    
    wire n1627, n3117, n3118, n3119, n3120, n3214, n3215, n3216, 
        n3217, n3218, n3219, n3220, n3221, n3222, n12324, n3223, 
        n3224, n3225, n3226, n3227, n10976, n44, n12216, n6_adj_1338, 
        n3376, n10904, n3230, n3243, n3369, n10895, n12215, n3368, 
        n11111, n11110, n3228, n3362, n3229, n35, n12314, n38, 
        n3158, n3147, n3146, n3145, n3148, n3378, n10871, n12057, 
        n3157, n3156, n3155, n12312, n3154, n12311, SRAM_DATA_out_14, 
        n12309, n63_adj_1339, SRAM_DATA_out_15, n11109, n11238, n12304, 
        n11237, n11235, n11234, n5_adj_1340, LOGIC_CLOCK_enable_48, 
        n11232, n11231, n11229, n11228, n11226, n11225, n12299, 
        n11223, SRAM_DATA_out_12, n11115, SRAM_DATA_out_11, SRAM_DATA_out_10, 
        SRAM_DATA_out_9, SRAM_DATA_out_8, SRAM_DATA_out_7, SRAM_DATA_out_6, 
        SRAM_DATA_out_5, SRAM_DATA_out_4, SRAM_DATA_out_3, SRAM_DATA_out_2, 
        SRAM_DATA_out_1, SRAM_DATA_out_0, PIC_DATA_IN_out_15, PIC_DATA_IN_out_14, 
        PIC_DATA_IN_out_13, PIC_DATA_IN_out_12, n11324, PIC_DATA_IN_out_11, 
        PIC_DATA_IN_out_10, PIC_DATA_IN_out_9, PIC_DATA_IN_out_8, PIC_DATA_IN_out_7, 
        PIC_DATA_IN_out_6, PIC_DATA_IN_out_5, PIC_DATA_IN_out_4, PIC_DATA_IN_out_3, 
        PIC_DATA_IN_out_2, PIC_DATA_IN_out_1, PIC_DATA_IN_out_0, n11122, 
        n11129, n11136, n11143, LOGIC_CLOCK_enable_168, n11150, n11157, 
        n11164, n11171, n12292, n11218, n11217, n11216, n11215, 
        n11213, n11212, n11210, n12291, n12290, n11209, n11207, 
        n12289, n12288, n11104, n11202, n11201, n11103, n11200, 
        n11199, n12287, n11197, n11102, n11196, n11194, BUS_ADDR_INTERNAL_18_derived_1, 
        n12284, n9991, n11189, n11188, n9990, n11187, n11186, 
        n11184, n11183, n11181, n11180, n11178, n11177, n11175, 
        n11174, n9989, n11172, n11758, LOGIC_CLOCK_enable_49, n9988, 
        n12280, n12279, n12278, n12277, n12276, n11167, n9987, 
        n11166, n11165, n11097, n12274, n11160, n11096, n11095, 
        n12273, n12272, n11094, n11159, n11158, n4_adj_1341, n11076, 
        n12271, n12270, n12269, n9986, n12268, n5_adj_1342, n12214, 
        n12213, n9985, n69, n12265, n12264, n12263, n12262, n12261, 
        n12259, n12258, n13160, n12253, n11066, n12252, n12251, 
        n12250, n12212, n12248, n12247, n12244, n100, n9924, n11485, 
        n12354, n12352, n12231, LOGIC_CLOCK_enable_26, n12227, n12223, 
        n12222, n12221, n12220;
    
    VHI i2 (.Z(VCC_net));
    BB SRAM_DATA_pad_12 (.I(BUS_data[12]), .T(SRAM_WE_c), .B(SRAM_DATA[12]), 
       .O(SRAM_DATA_out_12));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    CCU2D sub_676_add_2_7 (.A0(currPWMCount[5]), .B0(currPWMCountMax[5]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[6]), .B1(currPWMCountMax[6]), 
          .C1(GND_net), .D1(GND_net), .CIN(n9987), .COUT(n9988));
    defparam sub_676_add_2_7.INIT0 = 16'h5999;
    defparam sub_676_add_2_7.INIT1 = 16'h5999;
    defparam sub_676_add_2_7.INJECT1_0 = "NO";
    defparam sub_676_add_2_7.INJECT1_1 = "NO";
    LUT4 SRAM_WE_N_705_I_0_264_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(BUS_ADDR_INTERNAL_18_derived_1), .C(n12279), .D(n13140), .Z(lastAddress_31__N_788)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_264_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5c4;
    LUT4 lastAddress_i1_i1_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(lastAddress[0]), .D(n12277), .Z(n64)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i1_3_lut_3_lut_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i8230_3_lut_4_lut_4_lut (.A(n12344), .B(n3113), .C(n3129), .D(n12289), 
         .Z(n11122)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8230_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8273_3_lut_4_lut_4_lut (.A(n12344), .B(n3154), .C(n3170), .D(n12289), 
         .Z(n11165)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8273_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8203_3_lut_4_lut_4_lut (.A(n12344), .B(n3142), .C(n3158), .D(n12289), 
         .Z(n11095)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8203_3_lut_4_lut_4_lut.init = 16'hf0d8;
    SRAM RAM (.lastAddress({Open_0, lastAddress[30:17], Open_1, lastAddress[15], 
         Open_2, Open_3, Open_4, Open_5, Open_6, lastAddress[9:0]}), 
         .LOGIC_CLOCK(LOGIC_CLOCK), .lastAddress_31__N_872(lastAddress_31__N_872), 
         .n66({Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, 
         Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, 
         Open_20, Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
         Open_27, Open_28, Open_29, Open_30, Open_31, Open_32, n59, 
         n60, Open_33, Open_34, Open_35, Open_36}), .SRAM_OE_c(SRAM_OE_c), 
         .SRAM_WE_c(SRAM_WE_c), .lastAddress_31__N_785(lastAddress_31__N_785), 
         .lastAddress_31__N_845(lastAddress_31__N_845), .lastAddress_31__N_857(lastAddress_31__N_857), 
         .n55(n55), .lastAddress_31__N_786(lastAddress_31__N_786), .lastAddress_31__N_781(lastAddress_31__N_781), 
         .lastAddress_31__N_777(lastAddress_31__N_777), .BUS_DATA_INTERNAL({Open_37, 
         Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, Open_44, 
         Open_45, Open_46, Open_47, Open_48, BUS_DATA_INTERNAL_adj_1362[3:0]}), 
         .SRAM_DATA_out_0(SRAM_DATA_out_0), .SRAM_ADDR_c_0(SRAM_ADDR_c_0), 
         .n12269(n12269), .lastAddress_31__N_789(lastAddress_31__N_789), 
         .lastAddress_31__N_881(lastAddress_31__N_881), .n13160(n13160), 
         .lastAddress_31__N_875(lastAddress_31__N_875), .n61(n61), .lastAddress_31__N_860(lastAddress_31__N_860), 
         .n56(n56), .n12057(n12057), .SRAM_WE_N_704(SRAM_WE_N_704), .lastAddress_31__N_782(lastAddress_31__N_782), 
         .lastAddress_31__N_827(lastAddress_31__N_827), .n33(n33), .lastAddress_31__N_836(lastAddress_31__N_836), 
         .n48(n48), .BUS_DONE_INTERNAL(BUS_DONE_INTERNAL), .lastAddress_31__N_787(lastAddress_31__N_787), 
         .GND_net(GND_net), .lastAddress_31__N_884(lastAddress_31__N_884), 
         .n64(n64), .n39(n39), .n38(n38), .n35(n35), .n37(n37), .n36(n36), 
         .lastAddress_31__N_851(lastAddress_31__N_851), .lastAddress_31__N_779(lastAddress_31__N_779), 
         .lastAddress_31__N_774(lastAddress_31__N_774), .lastAddress_31__N_848(lastAddress_31__N_848), 
         .n52(n52), .lastAddress_31__N_778(lastAddress_31__N_778), .lastAddress_31__N_863(lastAddress_31__N_863), 
         .n57(n57), .lastAddress_31__N_783(lastAddress_31__N_783), .n42(n42), 
         .n41(n41), .n34(n34), .lastAddress_31__N_760(lastAddress_31__N_760), 
         .n43(n43), .n40(n40), .lastAddress_31__N_830(lastAddress_31__N_830), 
         .n46(n46), .\BUS_ADDR_INTERNAL[18]_derived_1 (BUS_ADDR_INTERNAL_18_derived_1), 
         .lastAddress_31__N_833(lastAddress_31__N_833), .n47(n47), .n44(n44), 
         .n45(n45), .lastAddress_31__N_790(lastAddress_31__N_790), .lastAddress_31__N_866(lastAddress_31__N_866), 
         .n58(n58), .n13141(n13141), .n87(n87), .\PWMArray[0][12] (\PWMArray[0] [12]), 
         .n12221(n12221), .\MATRIX_data[3] (MATRIX_data[3]), .lastAddress_31__N_784(lastAddress_31__N_784), 
         .\PWMArray[0][11] (\PWMArray[0] [11]), .\MATRIX_data[2] (MATRIX_data[2]), 
         .lastAddress_31__N_839(lastAddress_31__N_839), .n49(n49), .n12265(n12265), 
         .n12309(n12309), .SRAM_DATA_out_1(SRAM_DATA_out_1), .SRAM_DATA_out_2(SRAM_DATA_out_2), 
         .SRAM_DATA_out_3(SRAM_DATA_out_3), .SRAM_DATA_out_4(SRAM_DATA_out_4), 
         .SRAM_DATA_out_5(SRAM_DATA_out_5), .SRAM_DATA_out_6(SRAM_DATA_out_6), 
         .SRAM_DATA_out_7(SRAM_DATA_out_7), .\BUS_DATA_INTERNAL[8] (BUS_DATA_INTERNAL_adj_1362[8]), 
         .SRAM_DATA_out_8(SRAM_DATA_out_8), .\BUS_DATA_INTERNAL[9] (BUS_DATA_INTERNAL_adj_1362[9]), 
         .SRAM_DATA_out_9(SRAM_DATA_out_9), .\BUS_DATA_INTERNAL[10] (BUS_DATA_INTERNAL_adj_1362[10]), 
         .SRAM_DATA_out_10(SRAM_DATA_out_10), .\BUS_DATA_INTERNAL[11] (BUS_DATA_INTERNAL_adj_1362[11]), 
         .SRAM_DATA_out_11(SRAM_DATA_out_11), .\BUS_DATA_INTERNAL[12] (BUS_DATA_INTERNAL_adj_1362[12]), 
         .SRAM_DATA_out_12(SRAM_DATA_out_12), .\BUS_DATA_INTERNAL[13] (BUS_DATA_INTERNAL_adj_1362[13]), 
         .SRAM_DATA_out_13(SRAM_DATA_out_13), .\BUS_DATA_INTERNAL[14] (BUS_DATA_INTERNAL_adj_1362[14]), 
         .SRAM_DATA_out_14(SRAM_DATA_out_14), .\BUS_DATA_INTERNAL[15] (BUS_DATA_INTERNAL_adj_1362[15]), 
         .SRAM_DATA_out_15(SRAM_DATA_out_15), .SRAM_ADDR_c_1(SRAM_ADDR_c_1), 
         .SRAM_ADDR_c_2(SRAM_ADDR_c_2), .n12253(n12253), .SRAM_ADDR_c_3(SRAM_ADDR_c_3), 
         .n12264(n12264), .SRAM_ADDR_c_4(SRAM_ADDR_c_4), .n12259(n12259), 
         .SRAM_ADDR_c_5(SRAM_ADDR_c_5), .n12247(n12247), .SRAM_ADDR_c_6(SRAM_ADDR_c_6), 
         .n12252(n12252), .SRAM_ADDR_c_7(SRAM_ADDR_c_7), .n12263(n12263), 
         .SRAM_ADDR_c_8(SRAM_ADDR_c_8), .n12250(n12250), .SRAM_ADDR_c_9(SRAM_ADDR_c_9), 
         .n12271(n12271), .SRAM_ADDR_c_10(SRAM_ADDR_c_10), .n12268(n12268), 
         .SRAM_ADDR_c_11(SRAM_ADDR_c_11), .\BUS_addr[11] (BUS_addr[11]), 
         .SRAM_ADDR_c_12(SRAM_ADDR_c_12), .n12251(n12251), .SRAM_ADDR_c_13(SRAM_ADDR_c_13), 
         .\BUS_addr[13] (BUS_addr[13]), .SRAM_ADDR_c_14(SRAM_ADDR_c_14), 
         .\BUS_addr[14] (BUS_addr[14]), .SRAM_ADDR_c_15(SRAM_ADDR_c_15), 
         .n12270(n12270), .SRAM_ADDR_c_16(SRAM_ADDR_c_16), .n12262(n12262), 
         .SRAM_ADDR_c_17(SRAM_ADDR_c_17), .n12329(n12329), .\PWMArray[0][10] (\PWMArray[0] [10]), 
         .\MATRIX_data[1] (MATRIX_data[1]), .lastAddress_31__N_788(lastAddress_31__N_788), 
         .lastAddress_31__N_878(lastAddress_31__N_878), .lastAddress_31__N_869(lastAddress_31__N_869), 
         .lastAddress_31__N_780(lastAddress_31__N_780), .lastAddress_31__N_854(lastAddress_31__N_854), 
         .lastAddress_31__N_776(lastAddress_31__N_776), .lastAddress_31__N_842(lastAddress_31__N_842), 
         .lastAddress_31__N_775(lastAddress_31__N_775), .lastAddress_31__N_773(lastAddress_31__N_773), 
         .BUS_DIRECTION_INTERNAL(BUS_DIRECTION_INTERNAL), .\BUS_currGrantID[0] (BUS_currGrantID[0]), 
         .\BUS_currGrantID[1] (BUS_currGrantID[1]), .n12223(n12223), .n12217(n12217), 
         .n12216(n12216), .n54(n54), .MDM_done(MDM_done), .n1886(n1886), 
         .BUS_VALID_N_113(BUS_VALID_N_113), .n7(n7), .n63(n63_adj_1339), 
         .n12227(n12227), .LOGIC_CLOCK_enable_26(LOGIC_CLOCK_enable_26), 
         .LOGIC_CLOCK_enable_49(LOGIC_CLOCK_enable_49), .n12219(n12219), 
         .n1184(n1184), .LOGIC_CLOCK_enable_71(LOGIC_CLOCK_enable_71), .\lastAddress[12] (lastAddress[12]), 
         .\lastAddress[10] (lastAddress[10]), .n62(n62), .n12354(n12354), 
         .n63_adj_36(n63), .PWMArray_0__12__N_110(PWMArray_0__12__N_110), 
         .\lastAddress[16] (lastAddress[16]), .n2198(n2198), .BUS_VALID_N_1118(BUS_VALID_N_1118), 
         .n12220(n12220), .n4(n4), .\BUS_data[7] (BUS_data[7]), .n4_adj_37(n4_adj_1313), 
         .\BUS_data[6] (BUS_data[6]), .n4_adj_38(n4_adj_1314), .\BUS_data[5] (BUS_data[5]), 
         .n4_adj_39(n4_adj_1341), .\BUS_data[4] (BUS_data[4]), .transferMode_3__N_1115(transferMode_3__N_1115), 
         .\lastAddress[31] (lastAddress[31]), .n12258(n12258), .\PWMArray[0][9] (\PWMArray[0] [9]), 
         .\MATRIX_data[0] (MATRIX_data[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(192[7:23])
    LUT4 mux_531_i4_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[3]), .C(yOffset[3]), 
         .D(n12277), .Z(n2263)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i4_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i11_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(lastAddress[10]), .D(n12274), .Z(n54)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i11_3_lut_3_lut_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i8343_3_lut_4_lut_4_lut (.A(n12344), .B(n3362), .C(n3378), .D(n12289), 
         .Z(n11235)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8343_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8272_3_lut_4_lut_4_lut (.A(n12344), .B(n3119), .C(n3135), .D(n12289), 
         .Z(n11164)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8272_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8310_3_lut_4_lut_4_lut (.A(n12344), .B(n3250), .C(n3266), .D(n12289), 
         .Z(n11202)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8310_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), .B(n12280), 
         .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_836)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h2220;
    BB SRAM_DATA_pad_13 (.I(BUS_data[13]), .T(SRAM_WE_c), .B(SRAM_DATA[13]), 
       .O(SRAM_DATA_out_13));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i8339_3_lut_4_lut_4_lut (.A(n12344), .B(n3325), .C(n3341), .D(n12289), 
         .Z(n11231)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8339_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_193 (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n12273), .D(n13140), .Z(lastAddress_31__N_782)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+(D))) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_193.init = 16'hf5c4;
    LUT4 i8283_3_lut_4_lut_4_lut (.A(n12344), .B(n3364), .C(n3380), .D(n12289), 
         .Z(n11175)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8283_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3DX BUS_currGrantID__i1 (.D(BUS_currGrantID_3__N_72[0]), .SP(LOGIC_CLOCK_enable_168), 
            .CK(LOGIC_CLOCK), .CD(BUS_currGrantID_3__N_54), .Q(BUS_currGrantID[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam BUS_currGrantID__i1.GSR = "DISABLED";
    BB SRAM_DATA_pad_14 (.I(BUS_data[14]), .T(SRAM_WE_c), .B(SRAM_DATA[14]), 
       .O(SRAM_DATA_out_14));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    FD1P3DX BUS_DONE_OVERRIDE_38 (.D(n13160), .SP(LOGIC_CLOCK_enable_48), 
            .CK(LOGIC_CLOCK), .CD(BUS_currGrantID_3__N_54), .Q(BUS_DONE_OVERRIDE)) /* synthesis lse_init_val=0 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam BUS_DONE_OVERRIDE_38.GSR = "DISABLED";
    LUT4 i8294_3_lut_4_lut_4_lut (.A(n12344), .B(n3104), .C(n3120), .D(n12289), 
         .Z(n11186)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8294_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 SRAM_WE_N_705_I_0_256_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12274), .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_780)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_256_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hddd0;
    LUT4 lastAddress_i1_i16_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(lastAddress[15]), .D(n12290), .Z(n49)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i16_3_lut_3_lut_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i8226_3_lut_4_lut_4_lut (.A(n12344), .B(n3252), .C(n3268), .D(n12289), 
         .Z(n11118)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8226_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8291_3_lut_4_lut_4_lut (.A(n12344), .B(n3316), .C(n3332), .D(n12289), 
         .Z(n11183)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8291_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8279_3_lut_4_lut_4_lut (.A(n12344), .B(n3328), .C(n3344), .D(n12289), 
         .Z(n11171)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8279_3_lut_4_lut_4_lut.init = 16'hf0d8;
    BB SRAM_DATA_pad_15 (.I(BUS_data[15]), .T(SRAM_WE_c), .B(SRAM_DATA[15]), 
       .O(SRAM_DATA_out_15));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    CCU2D sub_676_add_2_3 (.A0(currPWMCount[1]), .B0(currPWMCountMax[1]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[2]), .B1(currPWMCountMax[2]), 
          .C1(GND_net), .D1(GND_net), .CIN(n9985), .COUT(n9986));
    defparam sub_676_add_2_3.INIT0 = 16'h5999;
    defparam sub_676_add_2_3.INIT1 = 16'h5999;
    defparam sub_676_add_2_3.INJECT1_0 = "NO";
    defparam sub_676_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_318 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .Z(n12344)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_318.init = 16'heeee;
    LUT4 i4705_2_lut_rep_218_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(n12289), .D(n12288), .Z(n12244)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4705_2_lut_rep_218_3_lut_4_lut.init = 16'hfff1;
    BB SRAM_DATA_pad_11 (.I(BUS_data[11]), .T(SRAM_WE_c), .B(SRAM_DATA[11]), 
       .O(SRAM_DATA_out_11));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    LUT4 i8320_3_lut_4_lut_4_lut (.A(n12344), .B(n3321), .C(n3337), .D(n12289), 
         .Z(n11212)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8320_3_lut_4_lut_4_lut.init = 16'hf0d8;
    BB SRAM_DATA_pad_10 (.I(BUS_data[10]), .T(SRAM_WE_c), .B(SRAM_DATA[10]), 
       .O(SRAM_DATA_out_10));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_9 (.I(BUS_data[9]), .T(SRAM_WE_c), .B(SRAM_DATA[9]), 
       .O(SRAM_DATA_out_9));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_8 (.I(BUS_data[8]), .T(SRAM_WE_c), .B(SRAM_DATA[8]), 
       .O(SRAM_DATA_out_8));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_7 (.I(BUS_data[7]), .T(SRAM_WE_c), .B(SRAM_DATA[7]), 
       .O(SRAM_DATA_out_7));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_6 (.I(BUS_data[6]), .T(SRAM_WE_c), .B(SRAM_DATA[6]), 
       .O(SRAM_DATA_out_6));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_5 (.I(BUS_data[5]), .T(SRAM_WE_c), .B(SRAM_DATA[5]), 
       .O(SRAM_DATA_out_5));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_4 (.I(BUS_data[4]), .T(SRAM_WE_c), .B(SRAM_DATA[4]), 
       .O(SRAM_DATA_out_4));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_3 (.I(BUS_data[3]), .T(SRAM_WE_c), .B(SRAM_DATA[3]), 
       .O(SRAM_DATA_out_3));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_2 (.I(BUS_data[2]), .T(SRAM_WE_c), .B(SRAM_DATA[2]), 
       .O(SRAM_DATA_out_2));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_1 (.I(BUS_data[1]), .T(SRAM_WE_c), .B(SRAM_DATA[1]), 
       .O(SRAM_DATA_out_1));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB SRAM_DATA_pad_0 (.I(BUS_data[0]), .T(SRAM_WE_c), .B(SRAM_DATA[0]), 
       .O(SRAM_DATA_out_0));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(52[2:11])
    BB PIC_DATA_IN_pad_15 (.I(BUS_data[15]), .T(PIC_OE_c), .B(PIC_DATA_IN[15]), 
       .O(PIC_DATA_IN_out_15));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_14 (.I(BUS_data[14]), .T(PIC_OE_c), .B(PIC_DATA_IN[14]), 
       .O(PIC_DATA_IN_out_14));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_13 (.I(BUS_data[13]), .T(PIC_OE_c), .B(PIC_DATA_IN[13]), 
       .O(PIC_DATA_IN_out_13));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_12 (.I(BUS_data[12]), .T(PIC_OE_c), .B(PIC_DATA_IN[12]), 
       .O(PIC_DATA_IN_out_12));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_11 (.I(BUS_data[11]), .T(PIC_OE_c), .B(PIC_DATA_IN[11]), 
       .O(PIC_DATA_IN_out_11));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_10 (.I(BUS_data[10]), .T(PIC_OE_c), .B(PIC_DATA_IN[10]), 
       .O(PIC_DATA_IN_out_10));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_9 (.I(BUS_data[9]), .T(PIC_OE_c), .B(PIC_DATA_IN[9]), 
       .O(PIC_DATA_IN_out_9));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_8 (.I(BUS_data[8]), .T(PIC_OE_c), .B(PIC_DATA_IN[8]), 
       .O(PIC_DATA_IN_out_8));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_7 (.I(BUS_data[7]), .T(PIC_OE_c), .B(PIC_DATA_IN[7]), 
       .O(PIC_DATA_IN_out_7));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_6 (.I(BUS_data[6]), .T(PIC_OE_c), .B(PIC_DATA_IN[6]), 
       .O(PIC_DATA_IN_out_6));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_5 (.I(BUS_data[5]), .T(PIC_OE_c), .B(PIC_DATA_IN[5]), 
       .O(PIC_DATA_IN_out_5));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_4 (.I(BUS_data[4]), .T(PIC_OE_c), .B(PIC_DATA_IN[4]), 
       .O(PIC_DATA_IN_out_4));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_3 (.I(BUS_data[3]), .T(PIC_OE_c), .B(PIC_DATA_IN[3]), 
       .O(PIC_DATA_IN_out_3));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_2 (.I(BUS_data[2]), .T(PIC_OE_c), .B(PIC_DATA_IN[2]), 
       .O(PIC_DATA_IN_out_2));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_1 (.I(BUS_data[1]), .T(PIC_OE_c), .B(PIC_DATA_IN[1]), 
       .O(PIC_DATA_IN_out_1));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    BB PIC_DATA_IN_pad_0 (.I(BUS_data[0]), .T(PIC_OE_c), .B(PIC_DATA_IN[0]), 
       .O(PIC_DATA_IN_out_0));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(97[2:13])
    OB UART_TX_pad (.I(GND_net), .O(UART_TX));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(11[3:10])
    OB Matrix_DATA_Out_pad_11 (.I(Matrix_DATA_Out_c_11), .O(Matrix_DATA_Out[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_10 (.I(Matrix_DATA_Out_c_10), .O(Matrix_DATA_Out[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_9 (.I(Matrix_DATA_Out_c_9), .O(Matrix_DATA_Out[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_8 (.I(Matrix_DATA_Out_c_8), .O(Matrix_DATA_Out[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_7 (.I(Matrix_DATA_Out_c_7), .O(Matrix_DATA_Out[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_6 (.I(Matrix_DATA_Out_c_6), .O(Matrix_DATA_Out[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_5 (.I(Matrix_DATA_Out_c_5), .O(Matrix_DATA_Out[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_4 (.I(Matrix_DATA_Out_c_4), .O(Matrix_DATA_Out[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_3 (.I(Matrix_DATA_Out_c_3), .O(Matrix_DATA_Out[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_2 (.I(Matrix_DATA_Out_c_2), .O(Matrix_DATA_Out[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_1 (.I(Matrix_DATA_Out_c_1), .O(Matrix_DATA_Out[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_DATA_Out_pad_0 (.I(Matrix_DATA_Out_c_0), .O(Matrix_DATA_Out[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(13[3:18])
    OB Matrix_LINE_SEL_Out_pad_3 (.I(GND_net), .O(Matrix_LINE_SEL_Out[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_LINE_SEL_Out_pad_2 (.I(Matrix_LINE_SEL_Out_c_2), .O(Matrix_LINE_SEL_Out[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_LINE_SEL_Out_pad_1 (.I(Matrix_LINE_SEL_Out_c_1), .O(Matrix_LINE_SEL_Out[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_LINE_SEL_Out_pad_0 (.I(Matrix_LINE_SEL_Out_c_0), .O(Matrix_LINE_SEL_Out[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(14[3:22])
    OB Matrix_CTRL_Out_pad_2 (.I(Matrix_CTRL_Out_c_2), .O(Matrix_CTRL_Out[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    OB Matrix_CTRL_Out_pad_1 (.I(Matrix_CTRL_Out_c_1), .O(Matrix_CTRL_Out[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    OB Matrix_CTRL_Out_pad_0 (.I(Matrix_CTRL_Out_c_0), .O(Matrix_CTRL_Out[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(15[3:18])
    OB SRAM_OE_pad (.I(SRAM_OE_c), .O(SRAM_OE));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(17[3:10])
    OB SRAM_WE_pad (.I(SRAM_WE_c), .O(SRAM_WE));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(18[3:10])
    OB SRAM_CE_pad (.I(GND_net), .O(SRAM_CE));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(19[3:10])
    OB SRAM_ADDR_pad_17 (.I(SRAM_ADDR_c_17), .O(SRAM_ADDR[17]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_16 (.I(SRAM_ADDR_c_16), .O(SRAM_ADDR[16]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_15 (.I(SRAM_ADDR_c_15), .O(SRAM_ADDR[15]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_14 (.I(SRAM_ADDR_c_14), .O(SRAM_ADDR[14]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_13 (.I(SRAM_ADDR_c_13), .O(SRAM_ADDR[13]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_12 (.I(SRAM_ADDR_c_12), .O(SRAM_ADDR[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_11 (.I(SRAM_ADDR_c_11), .O(SRAM_ADDR[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_10 (.I(SRAM_ADDR_c_10), .O(SRAM_ADDR[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_9 (.I(SRAM_ADDR_c_9), .O(SRAM_ADDR[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_8 (.I(SRAM_ADDR_c_8), .O(SRAM_ADDR[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_7 (.I(SRAM_ADDR_c_7), .O(SRAM_ADDR[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_6 (.I(SRAM_ADDR_c_6), .O(SRAM_ADDR[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_5 (.I(SRAM_ADDR_c_5), .O(SRAM_ADDR[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_4 (.I(SRAM_ADDR_c_4), .O(SRAM_ADDR[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_3 (.I(SRAM_ADDR_c_3), .O(SRAM_ADDR[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_2 (.I(SRAM_ADDR_c_2), .O(SRAM_ADDR[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_1 (.I(SRAM_ADDR_c_1), .O(SRAM_ADDR[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB SRAM_ADDR_pad_0 (.I(SRAM_ADDR_c_0), .O(SRAM_ADDR[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(21[3:12])
    OB PIC_READY_pad (.I(PIC_READY_c), .O(PIC_READY));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(28[3:12])
    OB LED_pad_7 (.I(GND_net), .O(LED[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_6 (.I(GND_net), .O(LED[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_5 (.I(GND_net), .O(LED[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_4 (.I(GND_net), .O(LED[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_3 (.I(GND_net), .O(LED[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_2 (.I(GND_net), .O(LED[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_1 (.I(GND_net), .O(LED[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    OB LED_pad_0 (.I(GND_net), .O(LED[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(30[3:6])
    IB CLK_pad (.I(CLK), .O(CLK_c));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    IB PIC_OE_pad (.I(PIC_OE), .O(PIC_OE_c));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(23[3:9])
    IB PIC_WE_IN_pad (.I(PIC_WE_IN), .O(PIC_WE_IN_c));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    IB PIC_ADDR_IN_pad_18 (.I(PIC_ADDR_IN[18]), .O(PIC_ADDR_IN_c_18));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_17 (.I(PIC_ADDR_IN[17]), .O(PIC_ADDR_IN_c_17));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_16 (.I(PIC_ADDR_IN[16]), .O(PIC_ADDR_IN_c_16));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_15 (.I(PIC_ADDR_IN[15]), .O(PIC_ADDR_IN_c_15));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_14 (.I(PIC_ADDR_IN[14]), .O(PIC_ADDR_IN_c_14));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_13 (.I(PIC_ADDR_IN[13]), .O(PIC_ADDR_IN_c_13));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_12 (.I(PIC_ADDR_IN[12]), .O(PIC_ADDR_IN_c_12));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_11 (.I(PIC_ADDR_IN[11]), .O(PIC_ADDR_IN_c_11));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_10 (.I(PIC_ADDR_IN[10]), .O(PIC_ADDR_IN_c_10));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_9 (.I(PIC_ADDR_IN[9]), .O(PIC_ADDR_IN_c_9));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_8 (.I(PIC_ADDR_IN[8]), .O(PIC_ADDR_IN_c_8));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_7 (.I(PIC_ADDR_IN[7]), .O(PIC_ADDR_IN_c_7));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_6 (.I(PIC_ADDR_IN[6]), .O(PIC_ADDR_IN_c_6));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_5 (.I(PIC_ADDR_IN[5]), .O(PIC_ADDR_IN_c_5));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_4 (.I(PIC_ADDR_IN[4]), .O(PIC_ADDR_IN_c_4));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_3 (.I(PIC_ADDR_IN[3]), .O(PIC_ADDR_IN_c_3));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_2 (.I(PIC_ADDR_IN[2]), .O(PIC_ADDR_IN_c_2));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_1 (.I(PIC_ADDR_IN[1]), .O(PIC_ADDR_IN_c_1));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    IB PIC_ADDR_IN_pad_0 (.I(PIC_ADDR_IN[0]), .O(PIC_ADDR_IN_c_0));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(26[3:14])
    LUT4 i8337_3_lut_4_lut_4_lut (.A(n12344), .B(n3361), .C(n3377), .D(n12289), 
         .Z(n11229)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8337_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i4754_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n2025), .D(n12279), .Z(GR_WR_ADDR[2])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A ((C)+!B))) */ ;
    defparam i4754_2_lut_3_lut_4_lut_4_lut.init = 16'h0c04;
    LUT4 i8289_3_lut_4_lut_4_lut (.A(n12344), .B(n3350), .C(n3366), .D(n12289), 
         .Z(n11181)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8289_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8219_3_lut_4_lut_4_lut (.A(n12344), .B(n3245), .C(n3261), .D(n12289), 
         .Z(n11111)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8219_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8132_1_lut_rep_283_2_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .Z(n12309)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i8132_1_lut_rep_283_2_lut.init = 16'h1111;
    LUT4 SRAM_WE_N_705_I_0_266_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12277), .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_790)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_266_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hddd0;
    GSR GSR_INST (.GSR(n12258));
    LUT4 i2_4_lut (.A(BUS_DATA_INTERNAL_adj_1362[13]), .B(MDM_data[13]), 
         .C(n12261), .D(PIC_data[13]), .Z(BUS_data[13])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut.init = 16'hffec;
    LUT4 i1_2_lut_4_lut (.A(n12265), .B(n12269), .C(n12218), .D(n4541), 
         .Z(n3278)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i8302_3_lut_4_lut_4_lut (.A(n12344), .B(n3352), .C(n3368), .D(n12289), 
         .Z(n11194)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8302_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8253_3_lut_4_lut_4_lut (.A(n12344), .B(n3221), .C(n3237), .D(n12289), 
         .Z(n11145)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8253_3_lut_4_lut_4_lut.init = 16'hf0d8;
    CCU2D sub_676_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n9991), .S0(n2589));
    defparam sub_676_add_2_cout.INIT0 = 16'h0000;
    defparam sub_676_add_2_cout.INIT1 = 16'h0000;
    defparam sub_676_add_2_cout.INJECT1_0 = "NO";
    defparam sub_676_add_2_cout.INJECT1_1 = "NO";
    LUT4 lastAddress_i1_i20_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[19]), 
         .Z(n45)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i20_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 SRAM_WE_N_705_I_0_236_2_lut_2_lut_3_lut_3_lut_4_lut_1_lut_1_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .Z(lastAddress_31__N_760)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam SRAM_WE_N_705_I_0_236_2_lut_2_lut_3_lut_3_lut_4_lut_1_lut_1_lut_4_lut.init = 16'h1111;
    LUT4 i1_2_lut_4_lut_adj_194 (.A(n12265), .B(n12269), .C(n12218), .D(n4537), 
         .Z(n3243)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam i1_2_lut_4_lut_adj_194.init = 16'h0400;
    LUT4 i2_4_lut_adj_195 (.A(BUS_DATA_INTERNAL_adj_1362[14]), .B(MDM_data[14]), 
         .C(n12261), .D(PIC_data[14]), .Z(BUS_data[14])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut_adj_195.init = 16'hffec;
    LUT4 i1_2_lut_4_lut_adj_196 (.A(n12265), .B(n12269), .C(n12218), .D(n4545), 
         .Z(n3277)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam i1_2_lut_4_lut_adj_196.init = 16'h0400;
    LUT4 i2_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DONE), .C(n12312), .D(n71), 
         .Z(n6)) /* synthesis lut_function=(!(A (C+!(D))+!A (B+(C+!(D))))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0b00;
    LUT4 i7268_2_lut_4_lut (.A(n13151), .B(BUS_ADDR_INTERNAL[16]), .C(n12332), 
         .D(n12290), .Z(n9924)) /* synthesis lut_function=(A (D)+!A !((C+!(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i7268_2_lut_4_lut.init = 16'hae00;
    CCU2D sub_676_add_2_13 (.A0(currPWMCount[11]), .B0(currPWMCountMax[11]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[12]), .B1(currPWMCountMax[12]), 
          .C1(GND_net), .D1(GND_net), .CIN(n9990), .COUT(n9991));
    defparam sub_676_add_2_13.INIT0 = 16'h5999;
    defparam sub_676_add_2_13.INIT1 = 16'h5999;
    defparam sub_676_add_2_13.INJECT1_0 = "NO";
    defparam sub_676_add_2_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_251_3_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[0]), .D(BUS_ADDR_INTERNAL_adj_1374[0]), .Z(n12277)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam i1_2_lut_rep_251_3_lut_4_lut_4_lut.init = 16'h6420;
    LUT4 i5_4_lut (.A(n69), .B(n7_adj_1308), .C(n10976), .D(n12253), 
         .Z(n10855)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i5_4_lut.init = 16'hfffe;
    CCU2D sub_676_add_2_11 (.A0(currPWMCount[9]), .B0(currPWMCountMax[9]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[10]), .B1(currPWMCountMax[10]), 
          .C1(GND_net), .D1(GND_net), .CIN(n9989), .COUT(n9990));
    defparam sub_676_add_2_11.INIT0 = 16'h5999;
    defparam sub_676_add_2_11.INIT1 = 16'h5999;
    defparam sub_676_add_2_11.INJECT1_0 = "NO";
    defparam sub_676_add_2_11.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_197 (.A(BUS_DATA_INTERNAL_adj_1362[8]), .B(MDM_data[8]), 
         .C(n12261), .D(PIC_data[8]), .Z(BUS_data[8])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut_adj_197.init = 16'hffec;
    CCU2D sub_676_add_2_9 (.A0(currPWMCount[7]), .B0(currPWMCountMax[7]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[8]), .B1(currPWMCountMax[8]), 
          .C1(GND_net), .D1(GND_net), .CIN(n9988), .COUT(n9989));
    defparam sub_676_add_2_9.INIT0 = 16'h5999;
    defparam sub_676_add_2_9.INIT1 = 16'h5999;
    defparam sub_676_add_2_9.INJECT1_0 = "NO";
    defparam sub_676_add_2_9.INJECT1_1 = "NO";
    LUT4 i4786_2_lut_rep_331 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[6]), .Z(n13146)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4786_2_lut_rep_331.init = 16'h2020;
    LUT4 i1_2_lut_rep_226_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[6]), .D(BUS_ADDR_INTERNAL[6]), 
         .Z(n12252)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_226_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4787_2_lut_rep_332 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[7]), .Z(n13147)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4787_2_lut_rep_332.init = 16'h2020;
    LUT4 i1_2_lut_rep_237_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[7]), .D(BUS_ADDR_INTERNAL[7]), .Z(n12263)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_237_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4783_2_lut_rep_333 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[3]), .Z(n13148)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4783_2_lut_rep_333.init = 16'h2020;
    LUT4 i2_4_lut_adj_198 (.A(BUS_DATA_INTERNAL_adj_1362[9]), .B(MDM_data[9]), 
         .C(n12261), .D(PIC_data[9]), .Z(BUS_data[9])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut_adj_198.init = 16'hffec;
    LUT4 i1_2_lut_rep_238_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[3]), .D(BUS_ADDR_INTERNAL[3]), .Z(n12264)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_238_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4781_2_lut_rep_334 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[1]), .Z(n13149)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4781_2_lut_rep_334.init = 16'h2020;
    LUT4 i4944_2_lut_rep_239_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[1]), .D(BUS_ADDR_INTERNAL[1]), .Z(n12265)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4944_2_lut_rep_239_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4795_2_lut_rep_335 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[15]), .Z(n13150)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4795_2_lut_rep_335.init = 16'h2020;
    LUT4 i4844_2_lut_rep_244_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[15]), .D(BUS_ADDR_INTERNAL[15]), 
         .Z(n12270)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4844_2_lut_rep_244_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4796_2_lut_rep_336 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[16]), .Z(n13151)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4796_2_lut_rep_336.init = 16'h2020;
    LUT4 i4845_2_lut_rep_236_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[16]), .D(BUS_ADDR_INTERNAL[16]), 
         .Z(n12262)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4845_2_lut_rep_236_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i2_4_lut_adj_199 (.A(BUS_DATA_INTERNAL_adj_1362[10]), .B(MDM_data[10]), 
         .C(n12261), .D(PIC_data[10]), .Z(BUS_data[10])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut_adj_199.init = 16'hffec;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DONE), .C(n12324), .D(state_adj_1377[4]), 
         .Z(n10904)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C)+!B (C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h040f;
    LUT4 i4782_2_lut_rep_337 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[2]), .Z(n13152)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4782_2_lut_rep_337.init = 16'h2020;
    LUT4 i2_2_lut_rep_227_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[2]), .D(BUS_ADDR_INTERNAL[2]), 
         .Z(n12253)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i2_2_lut_rep_227_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4784_2_lut_rep_338 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[4]), .Z(n13153)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4784_2_lut_rep_338.init = 16'h2020;
    LUT4 i1_2_lut_rep_233_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[4]), .D(BUS_ADDR_INTERNAL[4]), .Z(n12259)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_233_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4788_2_lut_rep_339 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[8]), .Z(n13154)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4788_2_lut_rep_339.init = 16'h2020;
    LUT4 i1_2_lut_rep_224_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[8]), .D(BUS_ADDR_INTERNAL[8]), 
         .Z(n12250)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_224_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4793_2_lut_3_lut_rep_340 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[13]), .Z(n13155)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4793_2_lut_3_lut_rep_340.init = 16'h2020;
    LUT4 i2_3_lut_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[13]), .D(BUS_ADDR_INTERNAL[13]), 
         .Z(BUS_addr[13])) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i2_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i8260_3_lut_4_lut_4_lut (.A(n12344), .B(n3222), .C(n3238), .D(n12289), 
         .Z(n11152)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8260_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i4791_2_lut_3_lut_rep_341 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[11]), .Z(n13156)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4791_2_lut_3_lut_rep_341.init = 16'h2020;
    LUT4 i2_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[11]), .D(BUS_ADDR_INTERNAL[11]), 
         .Z(BUS_addr[11])) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i2_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4794_2_lut_3_lut_rep_342 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[14]), .Z(n13157)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4794_2_lut_3_lut_rep_342.init = 16'h2020;
    LUT4 i2_4_lut_4_lut_4_lut_4_lut_adj_200 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[14]), .D(BUS_ADDR_INTERNAL[14]), 
         .Z(BUS_addr[14])) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i2_4_lut_4_lut_4_lut_4_lut_adj_200.init = 16'h7531;
    LUT4 i8210_3_lut_4_lut_4_lut (.A(n12344), .B(n3141), .C(n3157), .D(n12289), 
         .Z(n11102)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8210_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i2_4_lut_adj_201 (.A(BUS_DATA_INTERNAL_adj_1362[11]), .B(MDM_data[11]), 
         .C(n12261), .D(PIC_data[11]), .Z(BUS_data[11])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut_adj_201.init = 16'hffec;
    LUT4 i1_2_lut_rep_324 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(BUS_ADDR_INTERNAL[0]), .Z(n13139)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam i1_2_lut_rep_324.init = 16'h2020;
    LUT4 i1_2_lut_rep_243_3_lut_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(BUS_ADDR_INTERNAL[0]), .D(BUS_ADDR_INTERNAL_adj_1374[0]), 
         .Z(n12269)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam i1_2_lut_rep_243_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i1_2_lut_rep_325 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .C(reset), .Z(n13140)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam i1_2_lut_rep_325.init = 16'h2020;
    LUT4 i8682_2_lut_rep_232_2_lut_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(reset), .D(BUS_ADDR_INTERNAL_adj_1374[18]), 
         .Z(n12258)) /* synthesis lut_function=(A (B+!(C))+!A !((D)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam i8682_2_lut_rep_232_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h8ace;
    LUT4 i2_4_lut_adj_202 (.A(BUS_DATA_INTERNAL_adj_1362[12]), .B(MDM_data[12]), 
         .C(n12261), .D(PIC_data[12]), .Z(BUS_data[12])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i2_4_lut_adj_202.init = 16'hffec;
    LUT4 SRAM_WE_N_705_I_0_280_2_lut_2_lut_3_lut_3_lut_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(reset), .D(BUS_ADDR_INTERNAL_adj_1374[18]), 
         .Z(lastAddress_31__N_827)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam SRAM_WE_N_705_I_0_280_2_lut_2_lut_3_lut_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6420;
    LUT4 SRAM_WE_N_705_I_0_281_2_lut_3_lut_4_lut_4_lut_3_lut (.A(BUS_currGrantID[0]), 
         .B(BUS_currGrantID[1]), .C(reset), .Z(lastAddress_31__N_830)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam SRAM_WE_N_705_I_0_281_2_lut_3_lut_4_lut_4_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(n12288), .D(n12289), .Z(n4545)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i8621_3_lut_rep_326 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_DIRECTION_INTERNAL), .Z(n13141)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i8621_3_lut_rep_326.init = 16'h9b9b;
    LUT4 i4983_3_lut_4_lut_4_lut_then_2_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_DIRECTION_INTERNAL), .D(SRAM_WE_N_704), 
         .Z(n12354)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (B+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4983_3_lut_4_lut_4_lut_then_2_lut_4_lut.init = 16'h009b;
    LUT4 i1_2_lut_rep_235_3_lut_3_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_DIRECTION_INTERNAL), .D(BUS_ADDR_INTERNAL_adj_1374[18]), 
         .Z(n12261)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_235_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4464;
    LUT4 i4792_2_lut_rep_327 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[12]), .Z(n13142)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4792_2_lut_rep_327.init = 16'h2020;
    LUT4 i4841_2_lut_rep_225_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[12]), .D(BUS_ADDR_INTERNAL[12]), 
         .Z(n12251)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4841_2_lut_rep_225_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i3_4_lut (.A(n5), .B(BUS_DATA_INTERNAL_adj_1362[2]), .C(MATRIX_data[2]), 
         .D(n12261), .Z(BUS_data[2])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i3_4_lut.init = 16'hfefa;
    LUT4 i4790_2_lut_rep_328 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[10]), .Z(n13143)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4790_2_lut_rep_328.init = 16'h2020;
    LUT4 lastAddress_i1_i26_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[25]), 
         .Z(n39)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i26_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 i1_4_lut (.A(BUS_DATA_INTERNAL_adj_1373[2]), .B(n12215), .C(n12217), 
         .D(BUS_DATA_INTERNAL_adj_1354[2]), .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut.init = 16'heca0;
    FD1P3DX BUS_currGrantID__i2 (.D(BUS_currGrantID_3__N_72[1]), .SP(LOGIC_CLOCK_enable_168), 
            .CK(LOGIC_CLOCK), .CD(BUS_currGrantID_3__N_54), .Q(BUS_currGrantID[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam BUS_currGrantID__i2.GSR = "DISABLED";
    CCU2D sub_676_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(currPWMCount[0]), .B1(currPWMCountMax[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n9985));
    defparam sub_676_add_2_1.INIT0 = 16'h0000;
    defparam sub_676_add_2_1.INIT1 = 16'h5999;
    defparam sub_676_add_2_1.INJECT1_0 = "NO";
    defparam sub_676_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(n7167), .B(state_adj_1377[7]), .Z(state_7__N_1050[7])) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_242_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[10]), .D(BUS_ADDR_INTERNAL[10]), 
         .Z(n12268)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_242_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4789_2_lut_rep_329 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[9]), .Z(n13144)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4789_2_lut_rep_329.init = 16'h2020;
    LUT4 i1_2_lut_rep_245_4_lut_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_ADDR_INTERNAL_adj_1374[9]), .D(BUS_ADDR_INTERNAL[9]), 
         .Z(n12271)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_245_4_lut_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i1_2_lut_rep_222_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[9]), .D(BUS_ADDR_INTERNAL[9]), .Z(n12248)) /* synthesis lut_function=(A (B+!(C))+!A !((D)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_222_4_lut_4_lut_4_lut.init = 16'h8ace;
    LUT4 i1_2_lut_3_lut_4_lut_adj_203 (.A(n12344), .B(n12272), .C(n12273), 
         .D(n10895), .Z(n7_adj_1308)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i1_2_lut_3_lut_4_lut_adj_203.init = 16'hfdff;
    LUT4 lastAddress_i1_i6_3_lut_4_lut (.A(n12344), .B(n12272), .C(SRAM_WE_N_704), 
         .D(lastAddress[5]), .Z(n59)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam lastAddress_i1_i6_3_lut_4_lut.init = 16'hfd0d;
    LUT4 lastAddress_i1_i21_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[20]), 
         .Z(n44)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i21_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 i1_2_lut_3_lut_4_lut_3_lut_4_lut_adj_204 (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(n12288), .D(n12289), .Z(n4537)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_3_lut_4_lut_3_lut_4_lut_adj_204.init = 16'h0e00;
    LUT4 i4830_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(n12289), .D(n12288), .Z(n4541)) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4830_3_lut_3_lut_4_lut.init = 16'hf111;
    LUT4 lastAddress_i1_i25_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[24]), 
         .Z(n40)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i25_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i24_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[23]), 
         .Z(n41)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i24_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 i8266_3_lut_4_lut_4_lut (.A(n12344), .B(n3153), .C(n3169), .D(n12289), 
         .Z(n11158)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8266_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_4_lut_adj_205 (.A(n13147), .B(BUS_ADDR_INTERNAL[7]), .C(n12332), 
         .D(n12289), .Z(n69)) /* synthesis lut_function=(A+(B ((D)+!C)+!B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i1_2_lut_4_lut_adj_205.init = 16'hffae;
    LUT4 i1_2_lut_rep_322 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .Z(n12348)) /* synthesis lut_function=((B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_322.init = 16'hdddd;
    LUT4 i4619_2_lut_rep_288_3_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_DIRECTION_INTERNAL), .Z(n12314)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4619_2_lut_rep_288_3_lut.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_187_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(n71), .D(BUS_DONE), .Z(n12213)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_187_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i4607_2_lut_rep_273_3_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[0]), .Z(n12299)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4607_2_lut_rep_273_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_186_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(state_adj_1377[4]), .D(BUS_DONE), .Z(n12212)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_186_3_lut_4_lut.init = 16'h2f0f;
    LUT4 state_7__N_919_0__bdd_1_lut_3_lut_4_lut_3_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(BUS_DIRECTION_INTERNAL), .Z(n12057)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam state_7__N_919_0__bdd_1_lut_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 n23_bdd_2_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(state_adj_1377[1]), .D(BUS_DONE), .Z(n11758)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam n23_bdd_2_lut_3_lut_4_lut.init = 16'h0d0f;
    LUT4 i1_2_lut_rep_188_3_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_DONE), .Z(n12214)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_188_3_lut.init = 16'h2020;
    LUT4 i4785_2_lut_rep_330 (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[5]), .Z(n13145)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4785_2_lut_rep_330.init = 16'h2020;
    LUT4 i3050_1_lut (.A(BUS_currGrantID[1]), .Z(n5648)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i3050_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_221_4_lut_4_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[5]), .D(BUS_ADDR_INTERNAL[5]), .Z(n12247)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i1_2_lut_rep_221_4_lut_4_lut_4_lut.init = 16'h7531;
    LUT4 i4797_2_lut_rep_278_3_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[18]), .Z(n12304)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i4797_2_lut_rep_278_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_adj_206 (.A(n12215), .B(writeData[7]), .C(BUS_DATA_INTERNAL_adj_1354[7]), 
         .D(n12216), .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_206.init = 16'heca0;
    LUT4 i2343_2_lut_rep_260_3_lut_4_lut_3_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_ADDR_INTERNAL_adj_1374[18]), .Z(BUS_ADDR_INTERNAL_18_derived_1)) /* synthesis lut_function=(!(A (B+!(C))+!A (B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i2343_2_lut_rep_260_3_lut_4_lut_3_lut.init = 16'h3131;
    LUT4 i1_4_lut_adj_207 (.A(n12215), .B(writeData[6]), .C(BUS_DATA_INTERNAL_adj_1354[6]), 
         .D(n12216), .Z(n4_adj_1313)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_207.init = 16'heca0;
    LUT4 i1_4_lut_adj_208 (.A(n12215), .B(writeData[5]), .C(BUS_DATA_INTERNAL_adj_1354[5]), 
         .D(n12216), .Z(n4_adj_1314)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_208.init = 16'heca0;
    LUT4 i8239_3_lut_4_lut_4_lut (.A(n12344), .B(n3219), .C(n3235), .D(n12289), 
         .Z(n11131)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8239_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i4590_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n2025), .D(n12277), .Z(GR_WR_ADDR[0])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A ((C)+!B))) */ ;
    defparam i4590_2_lut_3_lut_4_lut_4_lut.init = 16'h0c04;
    LUT4 i8321_3_lut_4_lut_4_lut (.A(n12344), .B(n3356), .C(n3372), .D(n12289), 
         .Z(n11213)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8321_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8240_3_lut_4_lut_4_lut (.A(n12344), .B(n3254), .C(n3270), .D(n12289), 
         .Z(n11132)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8240_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i3_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(lastAddress[2]), .D(n12279), .Z(n62)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i3_3_lut_3_lut_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i8439_3_lut_4_lut_4_lut (.A(n12344), .B(n3108), .C(n3124), .D(n12289), 
         .Z(n11331)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8439_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8252_3_lut_4_lut_4_lut (.A(n12344), .B(n3151), .C(n3167), .D(n12289), 
         .Z(n11144)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8252_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_4_lut_adj_209 (.A(n12215), .B(writeData[4]), .C(BUS_DATA_INTERNAL_adj_1354[4]), 
         .D(n12216), .Z(n4_adj_1341)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_209.init = 16'heca0;
    LUT4 mux_531_i2_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[1]), .C(yOffset[1]), 
         .D(n12277), .Z(n2265)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i2_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i3_4_lut_adj_210 (.A(n5_adj_1307), .B(BUS_DATA_INTERNAL_adj_1362[1]), 
         .C(MATRIX_data[1]), .D(n12261), .Z(BUS_data[1])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i3_4_lut_adj_210.init = 16'hfefa;
    LUT4 i1_4_lut_adj_211 (.A(BUS_DATA_INTERNAL_adj_1373[1]), .B(n12215), 
         .C(n12217), .D(BUS_DATA_INTERNAL_adj_1354[1]), .Z(n5_adj_1307)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_211.init = 16'heca0;
    LUT4 mux_531_i5_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[4]), .C(yOffset[4]), 
         .D(n12277), .Z(n2262)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i5_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_212 (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n12279), .D(n13140), .Z(lastAddress_31__N_878)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_212.init = 16'h0a08;
    LUT4 i8265_3_lut_4_lut_4_lut (.A(n12344), .B(n3118), .C(n3134), .D(n12289), 
         .Z(n11157)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8265_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8305_3_lut_4_lut_4_lut (.A(n12344), .B(n3353), .C(n3369), .D(n12289), 
         .Z(n11197)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8305_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8232_3_lut_4_lut_4_lut (.A(n12344), .B(n3218), .C(n3234), .D(n12289), 
         .Z(n11124)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8232_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_531_i3_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[2]), .C(yOffset[2]), 
         .D(n12277), .Z(n2264)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i3_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8334_3_lut_4_lut_4_lut (.A(n12344), .B(n3358), .C(n3374), .D(n12289), 
         .Z(n11226)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8334_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i9_3_lut_4_lut_4_lut (.A(n12344), .B(lastAddress[8]), 
         .C(SRAM_WE_N_704), .D(n12273), .Z(n56)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam lastAddress_i1_i9_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i8275_3_lut_4_lut_4_lut (.A(n12344), .B(n3259), .C(n3275), .D(n12289), 
         .Z(n11167)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8275_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8209_3_lut_4_lut_4_lut (.A(n12344), .B(n3106), .C(n3122), .D(n12289), 
         .Z(n11101)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8209_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8433_3_lut_4_lut_4_lut (.A(n12344), .B(n3146), .C(n3162), .D(n12289), 
         .Z(n11325)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8433_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8435_3_lut_4_lut_4_lut (.A(n12344), .B(n3251), .C(n3267), .D(n12289), 
         .Z(n11327)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8435_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8218_3_lut_4_lut_4_lut (.A(n12344), .B(n3210), .C(n3226), .D(n12289), 
         .Z(n11110)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8218_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8288_3_lut_4_lut_4_lut (.A(n12344), .B(n3315), .C(n3331), .D(n12289), 
         .Z(n11180)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8288_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8282_3_lut_4_lut_4_lut (.A(n12344), .B(n3329), .C(n3345), .D(n12289), 
         .Z(n11174)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8282_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8317_3_lut_4_lut_4_lut (.A(n12344), .B(n3320), .C(n3336), .D(n12289), 
         .Z(n11209)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8317_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8325_3_lut_4_lut_4_lut (.A(n12344), .B(n3214), .C(n3230), .D(n12289), 
         .Z(n11217)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8325_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8202_3_lut_4_lut_4_lut (.A(n12344), .B(n3107), .C(n3123), .D(n12289), 
         .Z(n11094)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8202_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8224_3_lut_4_lut_4_lut (.A(n12344), .B(n3147), .C(n3163), .D(n12289), 
         .Z(n11116)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8224_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8297_3_lut_4_lut_4_lut (.A(n12344), .B(n3244), .C(n3260), .D(n12289), 
         .Z(n11189)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8297_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8233_3_lut_4_lut_4_lut (.A(n12344), .B(n3253), .C(n3269), .D(n12289), 
         .Z(n11125)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8233_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8258_3_lut_4_lut_4_lut (.A(n12344), .B(n3117), .C(n3133), .D(n12289), 
         .Z(n11150)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8258_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8212_3_lut_4_lut_4_lut (.A(n12344), .B(n3246), .C(n3262), .D(n12289), 
         .Z(n11104)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8212_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8268_3_lut_4_lut_4_lut (.A(n12344), .B(n3258), .C(n3274), .D(n12289), 
         .Z(n11160)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8268_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8309_3_lut_4_lut_4_lut (.A(n12344), .B(n3215), .C(n3231), .D(n12289), 
         .Z(n11201)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8309_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8345_3_lut_4_lut_4_lut (.A(n12344), .B(n3324), .C(n3340), .D(n12289), 
         .Z(n11237)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8345_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 SRAM_WE_N_705_I_0_250_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12280), .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_774)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_250_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hddd0;
    LUT4 i6_4_lut (.A(n13155), .B(n11066), .C(n12304), .D(n12344), .Z(n10871)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i6_4_lut.init = 16'h1000;
    LUT4 i8442_3_lut_4_lut_4_lut (.A(n12344), .B(n3248), .C(n3264), .D(n12289), 
         .Z(n11334)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8442_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8175_4_lut (.A(n13157), .B(n13156), .C(n12290), .D(n12280), 
         .Z(n11066)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8175_4_lut.init = 16'hfffe;
    LUT4 i8237_3_lut_4_lut_4_lut (.A(n12344), .B(n3114), .C(n3130), .D(n12289), 
         .Z(n11129)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8237_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8245_3_lut_4_lut_4_lut (.A(n12344), .B(n3150), .C(n3166), .D(n12289), 
         .Z(n11137)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8245_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8330_3_lut_4_lut_4_lut (.A(n12344), .B(n3322), .C(n3338), .D(n12289), 
         .Z(n11222)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8330_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8342_3_lut_4_lut_4_lut (.A(n12344), .B(n3327), .C(n3343), .D(n12289), 
         .Z(n11234)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8342_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 SRAM_WE_N_705_I_0_289_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12274), .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_854)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam SRAM_WE_N_705_I_0_289_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h2220;
    LUT4 i8292_3_lut_4_lut_4_lut (.A(n12344), .B(n3351), .C(n3367), .D(n12289), 
         .Z(n11184)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8292_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8441_3_lut_4_lut_4_lut (.A(n12344), .B(n3213), .C(n3229), .D(n12289), 
         .Z(n11333)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8441_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 SRAM_WE_N_705_I_0_284_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12290), .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_839)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam SRAM_WE_N_705_I_0_284_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h2220;
    LUT4 i8238_3_lut_4_lut_4_lut (.A(n12344), .B(n3149), .C(n3165), .D(n12289), 
         .Z(n11130)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8238_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8251_3_lut_4_lut_4_lut (.A(n12344), .B(n3116), .C(n3132), .D(n12289), 
         .Z(n11143)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8251_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n12344), .B(n10855), .C(n12292), .D(n12277), 
         .Z(n63_adj_1339)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffdf;
    LUT4 mux_531_i1_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[0]), .C(yOffset[0]), 
         .D(n12277), .Z(n2266)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i1_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8247_3_lut_4_lut_4_lut (.A(n12344), .B(n3255), .C(n3271), .D(n12289), 
         .Z(n11139)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8247_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i13_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(lastAddress[12]), .D(n12276), .Z(n52)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i13_3_lut_3_lut_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i8304_3_lut_4_lut_4_lut (.A(n12344), .B(n3318), .C(n3334), .D(n12289), 
         .Z(n11196)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8304_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8340_3_lut_4_lut_4_lut (.A(n12344), .B(n3360), .C(n3376), .D(n12289), 
         .Z(n11232)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8340_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8225_3_lut_4_lut_4_lut (.A(n12344), .B(n3217), .C(n3233), .D(n12289), 
         .Z(n11117)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8225_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8274_3_lut_4_lut_4_lut (.A(n12344), .B(n3224), .C(n3240), .D(n12289), 
         .Z(n11166)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8274_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8261_3_lut_4_lut_4_lut (.A(n12344), .B(n3257), .C(n3273), .D(n12289), 
         .Z(n11153)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8261_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_213 (.A(n12344), .B(n12291), 
         .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_781)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_213.init = 16'hddd0;
    LUT4 i8432_3_lut_4_lut_4_lut (.A(n12344), .B(n3111), .C(n3127), .D(n12289), 
         .Z(n11324)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8432_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8706_3_lut_4_lut_4_lut (.A(n12344), .B(n12304), .C(n1886), .D(BUS_VALID_N_113), 
         .Z(n11485)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;
    defparam i8706_3_lut_4_lut_4_lut.init = 16'h8088;
    LUT4 i8217_3_lut_4_lut_4_lut (.A(n12344), .B(n3140), .C(n3156), .D(n12289), 
         .Z(n11109)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8217_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8285_3_lut_4_lut_4_lut (.A(n12344), .B(n3314), .C(n3330), .D(n12289), 
         .Z(n11177)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8285_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8336_3_lut_4_lut_4_lut (.A(n12344), .B(n3326), .C(n3342), .D(n12289), 
         .Z(n11228)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8336_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8286_3_lut_4_lut_4_lut (.A(n12344), .B(n3349), .C(n3365), .D(n12289), 
         .Z(n11178)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8286_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8314_3_lut_4_lut_4_lut (.A(n12344), .B(n3319), .C(n3335), .D(n12289), 
         .Z(n11206)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8314_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8324_3_lut_4_lut_4_lut (.A(n12344), .B(n3144), .C(n3160), .D(n12289), 
         .Z(n11216)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8324_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_214 (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n12276), .D(n13140), .Z(lastAddress_31__N_848)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_214.init = 16'h0a08;
    LUT4 i8296_3_lut_4_lut_4_lut (.A(n12344), .B(n3209), .C(n3225), .D(n12289), 
         .Z(n11188)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8296_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_531_i7_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[6]), .C(yOffset[6]), 
         .D(n12277), .Z(n2260)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i7_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8205_3_lut_4_lut_4_lut (.A(n12344), .B(n3247), .C(n3263), .D(n12289), 
         .Z(n11097)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8205_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_rep_201_4_lut (.A(n12265), .B(n12277), .C(n10855), .D(n1184), 
         .Z(n12227)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam i1_2_lut_rep_201_4_lut.init = 16'hfb00;
    LUT4 i4758_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n2025), .D(n12289), .Z(GR_WR_ADDR[6])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A ((C)+!B))) */ ;
    defparam i4758_2_lut_3_lut_4_lut_4_lut.init = 16'h0c04;
    LUT4 i8295_3_lut_4_lut_4_lut (.A(n12344), .B(n3139), .C(n3155), .D(n12289), 
         .Z(n11187)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8295_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i7_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(lastAddress[6]), .D(n12289), .Z(n58)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i7_3_lut_3_lut_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i8204_3_lut_4_lut_4_lut (.A(n12344), .B(n3212), .C(n3228), .D(n12289), 
         .Z(n11096)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8204_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8323_3_lut_4_lut_4_lut (.A(n12344), .B(n3109), .C(n3125), .D(n12289), 
         .Z(n11215)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8323_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8315_3_lut_4_lut_4_lut (.A(n12344), .B(n3354), .C(n3370), .D(n12289), 
         .Z(n11207)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8315_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i3_4_lut_rep_205 (.A(n2589), .B(currPWMCount[13]), .C(currPWMCount[14]), 
         .D(currPWMCount[15]), .Z(n12231)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_rep_205.init = 16'hfffe;
    LUT4 i8307_3_lut_4_lut_4_lut (.A(n12344), .B(n3110), .C(n3126), .D(n12289), 
         .Z(n11199)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8307_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8434_3_lut_4_lut_4_lut (.A(n12344), .B(n3216), .C(n3232), .D(n12289), 
         .Z(n11326)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8434_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8216_3_lut_4_lut_4_lut (.A(n12344), .B(n3105), .C(n3121), .D(n12289), 
         .Z(n11108)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8216_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i17_3_lut_4_lut_4_lut (.A(n12344), .B(lastAddress[16]), 
         .C(SRAM_WE_N_704), .D(n12280), .Z(n48)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam lastAddress_i1_i17_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 SRAM_WE_N_705_I_0_251_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12290), .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_775)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_251_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hddd0;
    LUT4 mux_531_i8_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[7]), .C(yOffset[7]), 
         .D(n12277), .Z(n2259)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i8_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 SRAM_WE_N_705_I_0_260_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(BUS_ADDR_INTERNAL_18_derived_1), .C(n12289), .D(n13140), .Z(lastAddress_31__N_784)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_260_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5c4;
    LUT4 i8440_3_lut_4_lut_4_lut (.A(n12344), .B(n3143), .C(n3159), .D(n12289), 
         .Z(n11332)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8440_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8244_3_lut_4_lut_4_lut (.A(n12344), .B(n3115), .C(n3131), .D(n12289), 
         .Z(n11136)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8244_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8333_3_lut_4_lut_4_lut (.A(n12344), .B(n3323), .C(n3339), .D(n12289), 
         .Z(n11225)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8333_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8331_3_lut_4_lut_4_lut (.A(n12344), .B(n3357), .C(n3373), .D(n12289), 
         .Z(n11223)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8331_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8318_3_lut_4_lut_4_lut (.A(n12344), .B(n3355), .C(n3371), .D(n12289), 
         .Z(n11210)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8318_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8326_3_lut_4_lut_4_lut (.A(n12344), .B(n3249), .C(n3265), .D(n12289), 
         .Z(n11218)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8326_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8280_3_lut_4_lut_4_lut (.A(n12344), .B(n3363), .C(n3379), .D(n12289), 
         .Z(n11172)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8280_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_215 (.A(n12344), .B(n12277), 
         .C(BUS_ADDR_INTERNAL_18_derived_1), .D(n13140), .Z(lastAddress_31__N_884)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_215.init = 16'h2220;
    LUT4 i8223_3_lut_4_lut_4_lut (.A(n12344), .B(n3112), .C(n3128), .D(n12289), 
         .Z(n11115)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8223_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 lastAddress_i1_i10_3_lut_4_lut_4_lut (.A(n12344), .B(lastAddress[9]), 
         .C(SRAM_WE_N_704), .D(n12291), .Z(n55)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam lastAddress_i1_i10_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i8301_3_lut_4_lut_4_lut (.A(n12344), .B(n3317), .C(n3333), .D(n12289), 
         .Z(n11193)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8301_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8254_3_lut_4_lut_4_lut (.A(n12344), .B(n3256), .C(n3272), .D(n12289), 
         .Z(n11146)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8254_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8259_3_lut_4_lut_4_lut (.A(n12344), .B(n3152), .C(n3168), .D(n12289), 
         .Z(n11151)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8259_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_531_i6_3_lut_4_lut_4_lut (.A(n12344), .B(xOffset[5]), .C(yOffset[5]), 
         .D(n12277), .Z(n2261)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_531_i6_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8211_3_lut_4_lut_4_lut (.A(n12344), .B(n3211), .C(n3227), .D(n12289), 
         .Z(n11103)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8211_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8267_3_lut_4_lut_4_lut (.A(n12344), .B(n3223), .C(n3239), .D(n12289), 
         .Z(n11159)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8267_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8346_3_lut_4_lut_4_lut (.A(n12344), .B(n3359), .C(n3375), .D(n12289), 
         .Z(n11238)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8346_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_216 (.A(n12344), .B(BUS_ADDR_INTERNAL_18_derived_1), 
         .C(n12273), .D(n13140), .Z(lastAddress_31__N_860)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_216.init = 16'h0a08;
    LUT4 i8246_3_lut_4_lut_4_lut (.A(n12344), .B(n3220), .C(n3236), .D(n12289), 
         .Z(n11138)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8246_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i8308_3_lut_4_lut_4_lut (.A(n12344), .B(n3145), .C(n3161), .D(n12289), 
         .Z(n11200)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8308_3_lut_4_lut_4_lut.init = 16'hf0d8;
    CCU2D sub_676_add_2_5 (.A0(currPWMCount[3]), .B0(currPWMCountMax[3]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[4]), .B1(currPWMCountMax[4]), 
          .C1(GND_net), .D1(GND_net), .CIN(n9986), .COUT(n9987));
    defparam sub_676_add_2_5.INIT0 = 16'h5999;
    defparam sub_676_add_2_5.INIT1 = 16'h5999;
    defparam sub_676_add_2_5.INJECT1_0 = "NO";
    defparam sub_676_add_2_5.INJECT1_1 = "NO";
    LUT4 SRAM_WE_N_705_I_0_254_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(BUS_ADDR_INTERNAL_18_derived_1), .C(n12276), .D(n13140), .Z(lastAddress_31__N_778)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+(D))) */ ;
    defparam SRAM_WE_N_705_I_0_254_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5c4;
    LUT4 i8231_3_lut_4_lut_4_lut (.A(n12344), .B(n3148), .C(n3164), .D(n12289), 
         .Z(n11123)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam i8231_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 SRAM_WE_N_705_I_0_293_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(BUS_ADDR_INTERNAL_18_derived_1), .C(n12289), .D(n13140), .Z(lastAddress_31__N_866)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_705_I_0_293_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 i3_4_lut_adj_217 (.A(n5_adj_1340), .B(BUS_DATA_INTERNAL_adj_1362[0]), 
         .C(MATRIX_data[0]), .D(n12261), .Z(BUS_data[0])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i3_4_lut_adj_217.init = 16'hfefa;
    LUT4 i1_4_lut_adj_218 (.A(BUS_DATA_INTERNAL_adj_1373[0]), .B(n12215), 
         .C(n12217), .D(BUS_DATA_INTERNAL_adj_1354[0]), .Z(n5_adj_1340)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_218.init = 16'heca0;
    LUT4 i4_4_lut (.A(n12253), .B(n10976), .C(n12272), .D(n6_adj_1315), 
         .Z(n5045)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_219 (.A(n10871), .B(n13144), .C(n6_adj_1338), .D(n13158), 
         .Z(n10895)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i1_4_lut_adj_219.init = 16'h2000;
    LUT4 i2_4_lut_adj_220 (.A(n13142), .B(n11076), .C(n12274), .D(n12332), 
         .Z(n6_adj_1338)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[15:23])
    defparam i2_4_lut_adj_220.init = 16'h5010;
    LUT4 i8185_4_lut (.A(BUS_ADDR_INTERNAL[14]), .B(BUS_ADDR_INTERNAL[12]), 
         .C(BUS_ADDR_INTERNAL[9]), .D(n11004), .Z(n11076)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8185_4_lut.init = 16'hfffe;
    LUT4 i8117_2_lut (.A(BUS_ADDR_INTERNAL[11]), .B(BUS_ADDR_INTERNAL[13]), 
         .Z(n11004)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8117_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_221 (.A(n5_adj_1342), .B(BUS_DATA_INTERNAL_adj_1362[3]), 
         .C(MATRIX_data[3]), .D(n12261), .Z(BUS_data[3])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i3_4_lut_adj_221.init = 16'hfefa;
    LUT4 i1_4_lut_adj_222 (.A(BUS_DATA_INTERNAL_adj_1373[3]), .B(n12215), 
         .C(n12217), .D(BUS_DATA_INTERNAL_adj_1354[3]), .Z(n5_adj_1342)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(101[14:49])
    defparam i1_4_lut_adj_222.init = 16'heca0;
    LUT4 equal_781_i3_2_lut_rep_306 (.A(BUS_currGrantID[0]), .B(BUS_currGrantID[1]), 
         .Z(n12332)) /* synthesis lut_function=((B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(96[26:48])
    defparam equal_781_i3_2_lut_rep_306.init = 16'hdddd;
    LUT4 GR_WR_DOUT_9__I_0_i5_4_lut_4_lut (.A(n12265), .B(n1627), .C(n2262), 
         .D(GR_WR_DOUT[4]), .Z(otherData[4])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam GR_WR_DOUT_9__I_0_i5_4_lut_4_lut.init = 16'h7340;
    LUT4 GR_WR_DOUT_9__I_0_i6_4_lut_4_lut (.A(n12265), .B(n1627), .C(n2261), 
         .D(GR_WR_DOUT[5]), .Z(otherData[5])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam GR_WR_DOUT_9__I_0_i6_4_lut_4_lut.init = 16'h7340;
    LUT4 GR_WR_DOUT_9__I_0_i7_4_lut_4_lut (.A(n12265), .B(n1627), .C(n2260), 
         .D(GR_WR_DOUT[6]), .Z(otherData[6])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam GR_WR_DOUT_9__I_0_i7_4_lut_4_lut.init = 16'h7340;
    LUT4 GR_WR_DOUT_9__I_0_i8_4_lut_4_lut (.A(n12265), .B(n1627), .C(n2259), 
         .D(GR_WR_DOUT[7]), .Z(otherData[7])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam GR_WR_DOUT_9__I_0_i8_4_lut_4_lut.init = 16'h7340;
    PLL PLL_Ent (.LOGIC_CLOCK_N_116(LOGIC_CLOCK_N_116), .LOGIC_CLOCK(LOGIC_CLOCK), 
        .CLK_c(CLK_c), .PIXEL_CLOCK(PIXEL_CLOCK), .GND_net(GND_net), .PIXEL_CLOCK_N_302(PIXEL_CLOCK_N_302)) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(237[10:13])
    LUT4 lastAddress_i1_i30_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[29]), 
         .Z(n35)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i30_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i31_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[30]), 
         .Z(n34)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i31_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i28_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[27]), 
         .Z(n37)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i28_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i29_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[28]), 
         .Z(n36)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i29_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 i2_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(BUS_req[2]), .D(BUS_currGrantID_3__N_72[0]), .Z(LOGIC_CLOCK_enable_168)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 lastAddress_i1_i32_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), .B(BUS_currGrantID[0]), 
         .C(lastAddress[31]), .D(SRAM_WE_N_704), .Z(n33)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i32_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 lastAddress_i1_i27_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[26]), 
         .Z(n38)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i27_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i23_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[22]), 
         .Z(n42)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i23_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    LUT4 lastAddress_i1_i22_3_lut_3_lut_3_lut_4_lut (.A(BUS_currGrantID[1]), 
         .B(BUS_currGrantID[0]), .C(SRAM_WE_N_704), .D(lastAddress[21]), 
         .Z(n43)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(116[2] 134[9])
    defparam lastAddress_i1_i22_3_lut_3_lut_3_lut_4_lut.init = 16'hf101;
    MatrixBusHandler MDM (.\BUS_currGrantID[1] (BUS_currGrantID[1]), .\BUS_currGrantID[0] (BUS_currGrantID[0]), 
            .\BUS_ADDR_INTERNAL[13] (BUS_ADDR_INTERNAL[13]), .n13155(n13155), 
            .\BUS_ADDR_INTERNAL[14] (BUS_ADDR_INTERNAL[14]), .n13157(n13157), 
            .\BUS_ADDR_INTERNAL[11] (BUS_ADDR_INTERNAL[11]), .n13156(n13156), 
            .\BUS_ADDR_INTERNAL[12] (BUS_ADDR_INTERNAL[12]), .n13142(n13142), 
            .n12248(n12248), .n13158(n13158), .n12247(n12247), .n1627(n1627), 
            .GND_net(GND_net), .\BUS_ADDR_INTERNAL[10] (BUS_ADDR_INTERNAL[10]), 
            .n13143(n13143), .MATRIX_CURRROW({MATRIX_CURRROW}), .yOffset({yOffset}), 
            .n12342(n12342), .LOGIC_CLOCK(LOGIC_CLOCK), .n13160(n13160), 
            .LOGIC_CLOCK_enable_71(LOGIC_CLOCK_enable_71), .BUS_data({BUS_data}), 
            .\BUS_currGrantID_3__N_72[0] (BUS_currGrantID_3__N_72[0]), .\VRAM_ADDR[0] (VRAM_ADDR[0]), 
            .currReadRow({currReadRow}), .n12311(n12311), .n12284(n12284), 
            .n12253(n12253), .n12264(n12264), .n12259(n12259), .n3116(n3116), 
            .n3117(n3117), .n3118(n3118), .n3119(n3119), .n3112(n3112), 
            .n3113(n3113), .n3114(n3114), .n3115(n3115), .VRAM_WC(VRAM_WC), 
            .\BUS_ADDR_INTERNAL[0] (BUS_ADDR_INTERNAL[0]), .LOGIC_CLOCK_N_116(LOGIC_CLOCK_N_116), 
            .n12219(n12219), .n3132(n3132), .n3133(n3133), .n3134(n3134), 
            .n3135(n3135), .n3217(n3217), .n3218(n3218), .n3219(n3219), 
            .n3220(n3220), .n3322(n3322), .n3323(n3323), .n3324(n3324), 
            .n3325(n3325), .VRAM_DATA({VRAM_DATA}), .n12244(n12244), .n10871(n10871), 
            .n3167(n3167), .n3168(n3168), .n3169(n3169), .n3170(n3170), 
            .VCC_net(VCC_net), .n3027({n3027}), .\VRAM_ADDR[6] (VRAM_ADDR[6]), 
            .\VRAM_ADDR[5] (VRAM_ADDR[5]), .\VRAM_ADDR[4] (VRAM_ADDR[4]), 
            .MDM_done(MDM_done), .\VRAM_ADDR[3] (VRAM_ADDR[3]), .\VRAM_ADDR[2] (VRAM_ADDR[2]), 
            .xOffset({xOffset}), .\VRAM_ADDR[1] (VRAM_ADDR[1]), .n3035({n3035}), 
            .n3034({n3034}), .n3036({n3036}), .n3037({n3037}), .n3032({n3032}), 
            .n3031({n3031}), .n3033({n3033}), .n3029({n3029}), .n3028({n3028}), 
            .n3030({n3030}), .LOGIC_CLOCK_enable_26(LOGIC_CLOCK_enable_26), 
            .n5648(n5648), .\BUS_ADDR_INTERNAL[18] (BUS_ADDR_INTERNAL_adj_1374[18]), 
            .\BUS_ADDR_INTERNAL[16] (BUS_ADDR_INTERNAL_adj_1374[16]), .\BUS_ADDR_INTERNAL[16]_adj_19 (BUS_ADDR_INTERNAL[16]), 
            .\BUS_ADDR_INTERNAL[17] (BUS_ADDR_INTERNAL_adj_1374[17]), .\lastReadRow[3] (lastReadRow[3]), 
            .\lastReadRow[4] (lastReadRow[4]), .\BUS_ADDR_INTERNAL[15] (BUS_ADDR_INTERNAL[15]), 
            .\BUS_ADDR_INTERNAL[9] (BUS_ADDR_INTERNAL[9]), .\BUS_ADDR_INTERNAL[8] (BUS_ADDR_INTERNAL[8]), 
            .\BUS_ADDR_INTERNAL[7] (BUS_ADDR_INTERNAL[7]), .\BUS_ADDR_INTERNAL[6] (BUS_ADDR_INTERNAL[6]), 
            .\BUS_ADDR_INTERNAL[5] (BUS_ADDR_INTERNAL[5]), .\BUS_ADDR_INTERNAL[4] (BUS_ADDR_INTERNAL[4]), 
            .\BUS_ADDR_INTERNAL[3] (BUS_ADDR_INTERNAL[3]), .\BUS_ADDR_INTERNAL[2] (BUS_ADDR_INTERNAL[2]), 
            .\BUS_ADDR_INTERNAL[1] (BUS_ADDR_INTERNAL[1]), .\BUS_ADDR_INTERNAL[14]_adj_20 (BUS_ADDR_INTERNAL_adj_1374[14]), 
            .\BUS_ADDR_INTERNAL[15]_adj_21 (BUS_ADDR_INTERNAL_adj_1374[15]), 
            .\BUS_ADDR_INTERNAL[12]_adj_22 (BUS_ADDR_INTERNAL_adj_1374[12]), 
            .\BUS_ADDR_INTERNAL[13]_adj_23 (BUS_ADDR_INTERNAL_adj_1374[13]), 
            .\otherData[7] (otherData[7]), .\BUS_DATA_INTERNAL[7] (BUS_DATA_INTERNAL_adj_1354[7]), 
            .\otherData[6] (otherData[6]), .\BUS_DATA_INTERNAL[6] (BUS_DATA_INTERNAL_adj_1354[6]), 
            .\BUS_ADDR_INTERNAL[10]_adj_24 (BUS_ADDR_INTERNAL_adj_1374[10]), 
            .\BUS_ADDR_INTERNAL[11]_adj_25 (BUS_ADDR_INTERNAL_adj_1374[11]), 
            .\otherData[5] (otherData[5]), .\BUS_DATA_INTERNAL[5] (BUS_DATA_INTERNAL_adj_1354[5]), 
            .\BUS_ADDR_INTERNAL[8]_adj_26 (BUS_ADDR_INTERNAL_adj_1374[8]), 
            .\BUS_ADDR_INTERNAL[9]_adj_27 (BUS_ADDR_INTERNAL_adj_1374[9]), 
            .\otherData[4] (otherData[4]), .\BUS_DATA_INTERNAL[4] (BUS_DATA_INTERNAL_adj_1354[4]), 
            .\BUS_ADDR_INTERNAL[6]_adj_28 (BUS_ADDR_INTERNAL_adj_1374[6]), 
            .\BUS_ADDR_INTERNAL[7]_adj_29 (BUS_ADDR_INTERNAL_adj_1374[7]), 
            .\BUS_DATA_INTERNAL[3] (BUS_DATA_INTERNAL_adj_1354[3]), .n3365(n3365), 
            .n3366(n3366), .n3367(n3367), .n3368(n3368), .n3369(n3369), 
            .n3370(n3370), .n3371(n3371), .n3372(n3372), .n3373(n3373), 
            .n3374(n3374), .n3375(n3375), .n3376(n3376), .n3330(n3330), 
            .n3331(n3331), .n3332(n3332), .n3333(n3333), .n3334(n3334), 
            .n3335(n3335), .n3336(n3336), .n3337(n3337), .n3338(n3338), 
            .n3339(n3339), .n3340(n3340), .n3341(n3341), .n3349(n3349), 
            .n3350(n3350), .n3351(n3351), .n3352(n3352), .n3353(n3353), 
            .n3354(n3354), .n3355(n3355), .n3356(n3356), .n3357(n3357), 
            .n3358(n3358), .n3359(n3359), .n3360(n3360), .n3314(n3314), 
            .n3315(n3315), .n3316(n3316), .n3317(n3317), .n3318(n3318), 
            .n3319(n3319), .n3320(n3320), .n3321(n3321), .\BUS_DATA_INTERNAL[2] (BUS_DATA_INTERNAL_adj_1354[2]), 
            .n3361(n3361), .n3362(n3362), .n3363(n3363), .n3364(n3364), 
            .\BUS_DATA_INTERNAL[1] (BUS_DATA_INTERNAL_adj_1354[1]), .\BUS_ADDR_INTERNAL[4]_adj_30 (BUS_ADDR_INTERNAL_adj_1374[4]), 
            .\BUS_ADDR_INTERNAL[5]_adj_31 (BUS_ADDR_INTERNAL_adj_1374[5]), 
            .n3326(n3326), .n3327(n3327), .n3328(n3328), .n3329(n3329), 
            .n3342(n3342), .n3343(n3343), .n3344(n3344), .n3345(n3345), 
            .\BUS_ADDR_INTERNAL[2]_adj_32 (BUS_ADDR_INTERNAL_adj_1374[2]), 
            .\BUS_ADDR_INTERNAL[3]_adj_33 (BUS_ADDR_INTERNAL_adj_1374[3]), 
            .n3377(n3377), .n3378(n3378), .n3379(n3379), .n3380(n3380), 
            .n3260(n3260), .n3261(n3261), .n3262(n3262), .n3263(n3263), 
            .n3278(n3278), .n12277(n12277), .n12344(n12344), .n12292(n12292), 
            .\BUS_DATA_INTERNAL[0] (BUS_DATA_INTERNAL_adj_1354[0]), .n3264(n3264), 
            .n3265(n3265), .n3266(n3266), .n3267(n3267), .n3268(n3268), 
            .n3269(n3269), .n3270(n3270), .n3271(n3271), .n3225(n3225), 
            .n3226(n3226), .n3227(n3227), .n3228(n3228), .n3243(n3243), 
            .n3229(n3229), .n3230(n3230), .n3231(n3231), .n3232(n3232), 
            .n3233(n3233), .n3234(n3234), .n3235(n3235), .n3236(n3236), 
            .n3244(n3244), .n3245(n3245), .n3246(n3246), .n3247(n3247), 
            .n3277(n3277), .n3248(n3248), .n3249(n3249), .n3250(n3250), 
            .n3251(n3251), .n3252(n3252), .n3253(n3253), .n3254(n3254), 
            .n3255(n3255), .n3209(n3209), .n3210(n3210), .n3211(n3211), 
            .n3212(n3212), .n12269(n12269), .n3213(n3213), .n3214(n3214), 
            .n3215(n3215), .n3216(n3216), .n3256(n3256), .n3257(n3257), 
            .n3258(n3258), .n3259(n3259), .n3221(n3221), .n3222(n3222), 
            .n3223(n3223), .n3224(n3224), .n3237(n3237), .n3238(n3238), 
            .n3239(n3239), .n3240(n3240), .n3272(n3272), .n3273(n3273), 
            .n3274(n3274), .n3275(n3275), .n3155(n3155), .n3156(n3156), 
            .n3157(n3157), .n3158(n3158), .n3159(n3159), .n3160(n3160), 
            .n3161(n3161), .n3162(n3162), .n3163(n3163), .n3164(n3164), 
            .n3165(n3165), .n3166(n3166), .n3120(n3120), .n3121(n3121), 
            .n3122(n3122), .n3123(n3123), .n3124(n3124), .n3125(n3125), 
            .n3126(n3126), .n3127(n3127), .n3128(n3128), .n3129(n3129), 
            .n3130(n3130), .n3131(n3131), .n3139(n3139), .n3140(n3140), 
            .n3141(n3141), .n3142(n3142), .n3143(n3143), .n3144(n3144), 
            .n3145(n3145), .n3146(n3146), .n3147(n3147), .n3148(n3148), 
            .n3149(n3149), .n3150(n3150), .n3104(n3104), .n3105(n3105), 
            .n3106(n3106), .n3107(n3107), .n3108(n3108), .n3109(n3109), 
            .n3110(n3110), .n3111(n3111), .n3151(n3151), .n3152(n3152), 
            .n3153(n3153), .n3154(n3154), .n12309(n12309), .n13150(n13150), 
            .n13151(n13151), .reset(reset), .n13144(n13144), .n13154(n13154), 
            .LOGIC_CLOCK_enable_49(LOGIC_CLOCK_enable_49), .n11094(n11094), 
            .n11095(n11095), .n12263(n12263), .n11096(n11096), .n11097(n11097), 
            .n11150(n11150), .n11151(n11151), .n11152(n11152), .n11153(n11153), 
            .n11157(n11157), .n11158(n11158), .n11159(n11159), .n11160(n11160), 
            .n11164(n11164), .n11165(n11165), .n11166(n11166), .n11167(n11167), 
            .n1921(n1921), .n11171(n11171), .n11172(n11172), .n11174(n11174), 
            .n11175(n11175), .n11177(n11177), .n11178(n11178), .n11180(n11180), 
            .n11181(n11181), .n11183(n11183), .n11184(n11184), .n13146(n13146), 
            .n13147(n13147), .n13153(n13153), .n13145(n13145), .n13152(n13152), 
            .n13148(n13148), .n11101(n11101), .n11102(n11102), .n13139(n13139), 
            .n12299(n12299), .n11103(n11103), .n11104(n11104), .n12265(n12265), 
            .\MDM_data[13] (MDM_data[13]), .\MDM_data[14] (MDM_data[14]), 
            .n12261(n12261), .n100(n100), .\BUS_DATA_INTERNAL[15] (BUS_DATA_INTERNAL_adj_1362[15]), 
            .n12218(n12218), .n4537(n4537), .BUS_DONE(BUS_DONE), .n11186(n11186), 
            .n11187(n11187), .n4541(n4541), .n63(n63_adj_1339), .n1184(n1184), 
            .BUS_DONE_OUT_N_626(BUS_DONE_OUT_N_626), .n4545(n4545), .\MDM_data[8] (MDM_data[8]), 
            .n11188(n11188), .n11189(n11189), .\MDM_data[9] (MDM_data[9]), 
            .n11193(n11193), .n11194(n11194), .\MDM_data[10] (MDM_data[10]), 
            .n12329(n12329), .\MDM_data[11] (MDM_data[11]), .n13141(n13141), 
            .n12215(n12215), .n11196(n11196), .n11197(n11197), .n12332(n12332), 
            .n12352(n12352), .n12222(n12222), .n11199(n11199), .n11200(n11200), 
            .\BUS_ADDR_INTERNAL[18]_derived_1 (BUS_ADDR_INTERNAL_18_derived_1), 
            .\MDM_data[12] (MDM_data[12]), .n11201(n11201), .n11202(n11202), 
            .n11206(n11206), .n11207(n11207), .n11209(n11209), .n11210(n11210), 
            .n11212(n11212), .n11213(n11213), .n11215(n11215), .n11216(n11216), 
            .n11217(n11217), .n11218(n11218), .n12304(n12304), .\lastAddress[18] (lastAddress[18]), 
            .SRAM_WE_N_704(SRAM_WE_N_704), .n46(n46), .n2025(n2025), .n13140(n13140), 
            .lastAddress_31__N_789(lastAddress_31__N_789), .n12272(n12272), 
            .\BUS_addr[13] (BUS_addr[13]), .lastAddress_31__N_845(lastAddress_31__N_845), 
            .lastAddress_31__N_785(lastAddress_31__N_785), .n12288(n12288), 
            .lastAddress_31__N_863(lastAddress_31__N_863), .n12287(n12287), 
            .lastAddress_31__N_787(lastAddress_31__N_787), .lastAddress_31__N_783(lastAddress_31__N_783), 
            .n11222(n11222), .n11223(n11223), .\BUS_addr[11] (BUS_addr[11]), 
            .lastAddress_31__N_779(lastAddress_31__N_779), .lastAddress_31__N_851(lastAddress_31__N_851), 
            .lastAddress_31__N_869(lastAddress_31__N_869), .lastAddress_31__N_875(lastAddress_31__N_875), 
            .n12278(n12278), .lastAddress_31__N_881(lastAddress_31__N_881), 
            .lastAddress_31__N_777(lastAddress_31__N_777), .\BUS_addr[14] (BUS_addr[14]), 
            .lastAddress_31__N_842(lastAddress_31__N_842), .lastAddress_31__N_776(lastAddress_31__N_776), 
            .n12291(n12291), .lastAddress_31__N_857(lastAddress_31__N_857), 
            .lastAddress_31__N_872(lastAddress_31__N_872), .lastAddress_31__N_786(lastAddress_31__N_786), 
            .n11225(n11225), .n11226(n11226), .n11228(n11228), .n11229(n11229), 
            .n11231(n11231), .n11232(n11232), .n11234(n11234), .n11235(n11235), 
            .n11237(n11237), .n11238(n11238), .n11108(n11108), .n11109(n11109), 
            .n11110(n11110), .n11111(n11111), .n11115(n11115), .n11116(n11116), 
            .n12276(n12276), .n11012(n11012), .n12274(n12274), .n12273(n12273), 
            .n11117(n11117), .n11118(n11118), .n11122(n11122), .n11123(n11123), 
            .n10350(n10350), .n10349(n10349), .n11124(n11124), .n11125(n11125), 
            .n11129(n11129), .n11130(n11130), .n11131(n11131), .n11132(n11132), 
            .n12280(n12280), .n11324(n11324), .n11325(n11325), .n2266(n2266), 
            .n11326(n11326), .n11327(n11327), .n11136(n11136), .n11137(n11137), 
            .n10855(n10855), .\lastAddress[1] (lastAddress[1]), .n63_adj_34(n63), 
            .n2265(n2265), .n11331(n11331), .n11332(n11332), .n2264(n2264), 
            .n2263(n2263), .n11333(n11333), .n11334(n11334), .n11138(n11138), 
            .n11139(n11139), .n11143(n11143), .n11144(n11144), .n11145(n11145), 
            .n11146(n11146), .n12220(n12220), .WRITE_DONE(WRITE_DONE_adj_1337), 
            .WRITE_DONE_adj_35(WRITE_DONE), .n7(n7), .BUS_DONE_OVERRIDE(BUS_DONE_OVERRIDE), 
            .BUS_DONE_INTERNAL(BUS_DONE_INTERNAL), .\GR_WR_ADDR[6] (GR_WR_ADDR[6]), 
            .\GR_WR_ADDR[2] (GR_WR_ADDR[2]), .\GR_WR_ADDR[0] (GR_WR_ADDR[0]), 
            .\GR_WR_DOUT[7] (GR_WR_DOUT[7]), .\GR_WR_DOUT[6] (GR_WR_DOUT[6]), 
            .\GR_WR_DOUT[5] (GR_WR_DOUT[5]), .\GR_WR_DOUT[4] (GR_WR_DOUT[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    PIC PIC_BUS_INTERFACE (.GND_net(GND_net), .PIC_ADDR_IN_c_15(PIC_ADDR_IN_c_15), 
        .PIC_ADDR_IN_c_14(PIC_ADDR_IN_c_14), .PIC_ADDR_IN_c_13(PIC_ADDR_IN_c_13), 
        .PIC_ADDR_IN_c_12(PIC_ADDR_IN_c_12), .state({Open_49, Open_50, 
        Open_51, state_adj_1377[4], Open_52, Open_53, state_adj_1377[1], 
        Open_54}), .LOGIC_CLOCK(LOGIC_CLOCK), .\BUS_data[0] (BUS_data[0]), 
        .\BUS_ADDR_INTERNAL[0] (BUS_ADDR_INTERNAL_adj_1374[0]), .PIC_ADDR_IN_c_0(PIC_ADDR_IN_c_0), 
        .\BUS_req[2] (BUS_req[2]), .WRITE_DONE(WRITE_DONE_adj_1337), .transferMode_3__N_1115(transferMode_3__N_1115), 
        .n13160(n13160), .PIC_ADDR_IN_c_1(PIC_ADDR_IN_c_1), .PIC_ADDR_IN_c_2(PIC_ADDR_IN_c_2), 
        .PIC_ADDR_IN_c_3(PIC_ADDR_IN_c_3), .PIC_ADDR_IN_c_4(PIC_ADDR_IN_c_4), 
        .PIC_ADDR_IN_c_5(PIC_ADDR_IN_c_5), .PIC_ADDR_IN_c_6(PIC_ADDR_IN_c_6), 
        .PIC_ADDR_IN_c_7(PIC_ADDR_IN_c_7), .PIC_ADDR_IN_c_8(PIC_ADDR_IN_c_8), 
        .PIC_ADDR_IN_c_9(PIC_ADDR_IN_c_9), .PIC_ADDR_IN_c_10(PIC_ADDR_IN_c_10), 
        .PIC_ADDR_IN_c_11(PIC_ADDR_IN_c_11), .PIC_ADDR_IN_c_16(PIC_ADDR_IN_c_16), 
        .PIC_ADDR_IN_c_17(PIC_ADDR_IN_c_17), .PIC_ADDR_IN_c_18(PIC_ADDR_IN_c_18), 
        .n11758(n11758), .n5045(n5045), .n12252(n12252), .n12263(n12263), 
        .n87(n87), .BUS_VALID_N_1118(BUS_VALID_N_1118), .\BUS_currGrantID[0] (BUS_currGrantID[0]), 
        .\BUS_currGrantID[1] (BUS_currGrantID[1]), .n13158(n13158), .n12344(n12344), 
        .\BUS_ADDR_INTERNAL[18] (BUS_ADDR_INTERNAL_adj_1374[18]), .n12309(n12309), 
        .\BUS_ADDR_INTERNAL[15] (BUS_ADDR_INTERNAL[15]), .n13150(n13150), 
        .\BUS_ADDR_INTERNAL[16] (BUS_ADDR_INTERNAL[16]), .n13151(n13151), 
        .\BUS_ADDR_INTERNAL[13] (BUS_ADDR_INTERNAL[13]), .n13155(n13155), 
        .\BUS_ADDR_INTERNAL[14] (BUS_ADDR_INTERNAL[14]), .n13157(n13157), 
        .\BUS_ADDR_INTERNAL[11] (BUS_ADDR_INTERNAL[11]), .n13156(n13156), 
        .\BUS_ADDR_INTERNAL[12] (BUS_ADDR_INTERNAL[12]), .n13142(n13142), 
        .\BUS_ADDR_INTERNAL[9] (BUS_ADDR_INTERNAL[9]), .n13144(n13144), 
        .\BUS_ADDR_INTERNAL[10] (BUS_ADDR_INTERNAL[10]), .n13143(n13143), 
        .\BUS_ADDR_INTERNAL[8] (BUS_ADDR_INTERNAL[8]), .n13154(n13154), 
        .PIC_DATA_IN_out_15(PIC_DATA_IN_out_15), .PIC_DATA_IN_out_13(PIC_DATA_IN_out_13), 
        .PIC_DATA_IN_out_14(PIC_DATA_IN_out_14), .PIC_DATA_IN_out_11(PIC_DATA_IN_out_11), 
        .PIC_DATA_IN_out_12(PIC_DATA_IN_out_12), .PIC_DATA_IN_out_9(PIC_DATA_IN_out_9), 
        .PIC_DATA_IN_out_10(PIC_DATA_IN_out_10), .PIC_DATA_IN_out_8(PIC_DATA_IN_out_8), 
        .PIC_READY_c(PIC_READY_c), .BUS_DIRECTION_INTERNAL(BUS_DIRECTION_INTERNAL), 
        .n2198(n2198), .\BUS_data[1] (BUS_data[1]), .\BUS_data[2] (BUS_data[2]), 
        .\BUS_data[3] (BUS_data[3]), .\BUS_ADDR_INTERNAL[1] (BUS_ADDR_INTERNAL_adj_1374[1]), 
        .\BUS_ADDR_INTERNAL[2] (BUS_ADDR_INTERNAL_adj_1374[2]), .\BUS_ADDR_INTERNAL[3] (BUS_ADDR_INTERNAL_adj_1374[3]), 
        .\BUS_ADDR_INTERNAL[4] (BUS_ADDR_INTERNAL_adj_1374[4]), .\BUS_ADDR_INTERNAL[5] (BUS_ADDR_INTERNAL_adj_1374[5]), 
        .\BUS_ADDR_INTERNAL[6] (BUS_ADDR_INTERNAL_adj_1374[6]), .\BUS_ADDR_INTERNAL[7] (BUS_ADDR_INTERNAL_adj_1374[7]), 
        .\BUS_ADDR_INTERNAL[8]_adj_1 (BUS_ADDR_INTERNAL_adj_1374[8]), .\BUS_ADDR_INTERNAL[9]_adj_2 (BUS_ADDR_INTERNAL_adj_1374[9]), 
        .\BUS_ADDR_INTERNAL[10]_adj_3 (BUS_ADDR_INTERNAL_adj_1374[10]), .\BUS_ADDR_INTERNAL[11]_adj_4 (BUS_ADDR_INTERNAL_adj_1374[11]), 
        .\BUS_ADDR_INTERNAL[12]_adj_5 (BUS_ADDR_INTERNAL_adj_1374[12]), .\BUS_ADDR_INTERNAL[13]_adj_6 (BUS_ADDR_INTERNAL_adj_1374[13]), 
        .\BUS_ADDR_INTERNAL[14]_adj_7 (BUS_ADDR_INTERNAL_adj_1374[14]), .\BUS_ADDR_INTERNAL[15]_adj_8 (BUS_ADDR_INTERNAL_adj_1374[15]), 
        .\BUS_ADDR_INTERNAL[16]_adj_9 (BUS_ADDR_INTERNAL_adj_1374[16]), .\BUS_ADDR_INTERNAL[17] (BUS_ADDR_INTERNAL_adj_1374[17]), 
        .PIC_DATA_IN_out_3(PIC_DATA_IN_out_3), .PIC_WE_IN_c(PIC_WE_IN_c), 
        .PIC_DATA_IN_out_6(PIC_DATA_IN_out_6), .n12276(n12276), .n12274(n12274), 
        .n12291(n12291), .\BUS_ADDR_INTERNAL[5]_adj_10 (BUS_ADDR_INTERNAL[5]), 
        .n12272(n12272), .\BUS_ADDR_INTERNAL[6]_adj_11 (BUS_ADDR_INTERNAL[6]), 
        .n12289(n12289), .\BUS_ADDR_INTERNAL[7]_adj_12 (BUS_ADDR_INTERNAL[7]), 
        .n12288(n12288), .PIC_DATA_IN_out_5(PIC_DATA_IN_out_5), .PIC_DATA_IN_out_7(PIC_DATA_IN_out_7), 
        .\BUS_ADDR_INTERNAL[3]_adj_13 (BUS_ADDR_INTERNAL[3]), .n12287(n12287), 
        .n12290(n12290), .\BUS_data[4] (BUS_data[4]), .\BUS_data[5] (BUS_data[5]), 
        .\BUS_data[6] (BUS_data[6]), .\BUS_data[7] (BUS_data[7]), .\BUS_ADDR_INTERNAL[1]_adj_14 (BUS_ADDR_INTERNAL[1]), 
        .n12292(n12292), .\writeData[4] (writeData[4]), .\writeData[5] (writeData[5]), 
        .\writeData[6] (writeData[6]), .\writeData[7] (writeData[7]), .n12280(n12280), 
        .n1921(n1921), .n12222(n12222), .n2025(n2025), .LOGIC_CLOCK_enable_26(LOGIC_CLOCK_enable_26), 
        .\BUS_ADDR_INTERNAL[2]_adj_15 (BUS_ADDR_INTERNAL[2]), .n12279(n12279), 
        .\BUS_ADDR_INTERNAL[4]_adj_16 (BUS_ADDR_INTERNAL[4]), .n12278(n12278), 
        .n13147(n13147), .\state[7] (state_adj_1377[7]), .\state_7__N_1050[7] (state_7__N_1050[7]), 
        .n12273(n12273), .n13145(n13145), .n13146(n13146), .n13148(n13148), 
        .n13153(n13153), .n13149(n13149), .n13152(n13152), .\BUS_ADDR_INTERNAL[0]_adj_17 (BUS_ADDR_INTERNAL[0]), 
        .n12299(n12299), .PIC_DATA_IN_out_1(PIC_DATA_IN_out_1), .PIC_DATA_IN_out_2(PIC_DATA_IN_out_2), 
        .PIC_DATA_IN_out_4(PIC_DATA_IN_out_4), .n12223(n12223), .n13141(n13141), 
        .n11485(n11485), .n12219(n12219), .LOGIC_CLOCK_enable_48(LOGIC_CLOCK_enable_48), 
        .n7167(n7167), .n12213(n12213), .n12314(n12314), .\BUS_DATA_INTERNAL[2] (BUS_DATA_INTERNAL_adj_1373[2]), 
        .n6(n6), .\BUS_currGrantID_3__N_72[0] (BUS_currGrantID_3__N_72[0]), 
        .\BUS_currGrantID_3__N_72[1] (BUS_currGrantID_3__N_72[1]), .n12352(n12352), 
        .n71(n71), .PIC_OE_c(PIC_OE_c), .n12312(n12312), .n12214(n12214), 
        .n12324(n12324), .PIC_DATA_IN_out_0(PIC_DATA_IN_out_0), .n12212(n12212), 
        .n12348(n12348), .n13139(n13139), .n6_adj_18(n6_adj_1315), .\BUS_DATA_INTERNAL[1] (BUS_DATA_INTERNAL_adj_1373[1]), 
        .n10895(n10895), .n69(n69), .n1184(n1184), .BUS_currGrantID_3__N_54(BUS_currGrantID_3__N_54), 
        .BUS_DONE(BUS_DONE), .\BUS_DATA_INTERNAL[0] (BUS_DATA_INTERNAL_adj_1373[0]), 
        .n12250(n12250), .n12217(n12217), .\PIC_data[9] (PIC_data[9]), 
        .\PIC_data[11] (PIC_data[11]), .\PIC_data[10] (PIC_data[10]), .n100(n100), 
        .\PIC_data[12] (PIC_data[12]), .\PIC_data[8] (PIC_data[8]), .\PIC_data[13] (PIC_data[13]), 
        .\PIC_data[14] (PIC_data[14]), .SRAM_WE_N_704(SRAM_WE_N_704), .\lastAddress[4] (lastAddress[4]), 
        .n60(n60), .n10904(n10904), .\lastAddress[7] (lastAddress[7]), 
        .n57(n57), .\lastAddress[3] (lastAddress[3]), .n61(n61), .\lastAddress[17] (lastAddress[17]), 
        .n47(n47), .n13140(n13140), .n12304(n12304), .lastAddress_31__N_833(lastAddress_31__N_833), 
        .lastAddress_31__N_773(lastAddress_31__N_773), .n9924(n9924), .BUS_DONE_OUT_N_626(BUS_DONE_OUT_N_626), 
        .\BUS_DATA_INTERNAL[3] (BUS_DATA_INTERNAL_adj_1373[3]), .n12332(n12332), 
        .n10976(n10976), .n11012(n11012));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(211[21:36])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    MatrixDriver MD (.PIXEL_CLOCK(PIXEL_CLOCK), .\BUS_currGrantID[0] (BUS_currGrantID[0]), 
            .\BUS_currGrantID[1] (BUS_currGrantID[1]), .GND_net(GND_net), 
            .BUS_VALID_N_113(BUS_VALID_N_113), .Matrix_LINE_SEL_Out_c_0(Matrix_LINE_SEL_Out_c_0), 
            .\BUS_ADDR_INTERNAL[18] (BUS_ADDR_INTERNAL_adj_1374[18]), .n12309(n12309), 
            .Matrix_CTRL_Out_c_1(Matrix_CTRL_Out_c_1), .PIXEL_CLOCK_N_302(PIXEL_CLOCK_N_302), 
            .\BUS_ADDR_INTERNAL[16] (BUS_ADDR_INTERNAL[16]), .n13151(n13151), 
            .n13158(n13158), .n12344(n12344), .currPWMCount({currPWMCount}), 
            .LOGIC_CLOCK(LOGIC_CLOCK), .\BUS_ADDR_INTERNAL[14] (BUS_ADDR_INTERNAL[14]), 
            .n13157(n13157), .\BUS_ADDR_INTERNAL[15] (BUS_ADDR_INTERNAL[15]), 
            .n13150(n13150), .WRITE_DONE(WRITE_DONE), .LOGIC_CLOCK_N_116(LOGIC_CLOCK_N_116), 
            .PWMArray_0__12__N_110(PWMArray_0__12__N_110), .n13160(n13160), 
            .\PWMArray[0][12] (\PWMArray[0] [12]), .\BUS_data[3] (BUS_data[3]), 
            .\currPWMCountMax[0] (currPWMCountMax[0]), .\BUS_ADDR_INTERNAL[12] (BUS_ADDR_INTERNAL[12]), 
            .n13142(n13142), .\BUS_ADDR_INTERNAL[13] (BUS_ADDR_INTERNAL[13]), 
            .n13155(n13155), .\BUS_ADDR_INTERNAL[10] (BUS_ADDR_INTERNAL[10]), 
            .n13143(n13143), .\BUS_ADDR_INTERNAL[11] (BUS_ADDR_INTERNAL[11]), 
            .n13156(n13156), .\PWMArray[0][11] (\PWMArray[0] [11]), .\BUS_data[2] (BUS_data[2]), 
            .\BUS_ADDR_INTERNAL[8] (BUS_ADDR_INTERNAL[8]), .n13154(n13154), 
            .\BUS_ADDR_INTERNAL[9] (BUS_ADDR_INTERNAL[9]), .n13144(n13144), 
            .\BUS_ADDR_INTERNAL[7] (BUS_ADDR_INTERNAL[7]), .n13147(n13147), 
            .MATRIX_CURRROW({MATRIX_CURRROW}), .\PWMArray[0][9] (\PWMArray[0] [9]), 
            .\BUS_data[0] (BUS_data[0]), .\PWMArray[0][10] (\PWMArray[0] [10]), 
            .\BUS_data[1] (BUS_data[1]), .\currPWMCountMax[2] (currPWMCountMax[2]), 
            .\currPWMCountMax[5] (currPWMCountMax[5]), .\currPWMCountMax[1] (currPWMCountMax[1]), 
            .\currPWMCountMax[4] (currPWMCountMax[4]), .\currPWMCountMax[3] (currPWMCountMax[3]), 
            .\currPWMCountMax[6] (currPWMCountMax[6]), .Matrix_LINE_SEL_Out_c_1(Matrix_LINE_SEL_Out_c_1), 
            .n1886(n1886), .\currPWMCountMax[12] (currPWMCountMax[12]), 
            .Matrix_CTRL_Out_c_2(Matrix_CTRL_Out_c_2), .\currPWMCountMax[11] (currPWMCountMax[11]), 
            .\currPWMCountMax[10] (currPWMCountMax[10]), .\currPWMCountMax[9] (currPWMCountMax[9]), 
            .\currPWMCountMax[8] (currPWMCountMax[8]), .\currPWMCountMax[7] (currPWMCountMax[7]), 
            .\BUS_ADDR_INTERNAL[5] (BUS_ADDR_INTERNAL[5]), .n13145(n13145), 
            .\BUS_ADDR_INTERNAL[6] (BUS_ADDR_INTERNAL[6]), .n13146(n13146), 
            .\BUS_ADDR_INTERNAL[3] (BUS_ADDR_INTERNAL[3]), .n13148(n13148), 
            .\BUS_ADDR_INTERNAL[4] (BUS_ADDR_INTERNAL[4]), .n13153(n13153), 
            .\BUS_ADDR_INTERNAL[1] (BUS_ADDR_INTERNAL[1]), .n13149(n13149), 
            .\BUS_ADDR_INTERNAL[2] (BUS_ADDR_INTERNAL[2]), .n13152(n13152), 
            .\BUS_ADDR_INTERNAL[0] (BUS_ADDR_INTERNAL[0]), .n12299(n12299), 
            .currReadRow({currReadRow}), .n12231(n12231), .Matrix_DATA_Out_c_11(Matrix_DATA_Out_c_11), 
            .Matrix_DATA_Out_c_10(Matrix_DATA_Out_c_10), .Matrix_DATA_Out_c_9(Matrix_DATA_Out_c_9), 
            .Matrix_DATA_Out_c_8(Matrix_DATA_Out_c_8), .Matrix_DATA_Out_c_7(Matrix_DATA_Out_c_7), 
            .Matrix_DATA_Out_c_6(Matrix_DATA_Out_c_6), .Matrix_DATA_Out_c_5(Matrix_DATA_Out_c_5), 
            .Matrix_DATA_Out_c_4(Matrix_DATA_Out_c_4), .Matrix_DATA_Out_c_3(Matrix_DATA_Out_c_3), 
            .Matrix_DATA_Out_c_2(Matrix_DATA_Out_c_2), .Matrix_DATA_Out_c_1(Matrix_DATA_Out_c_1), 
            .Matrix_DATA_Out_c_0(Matrix_DATA_Out_c_0), .Matrix_LINE_SEL_Out_c_2(Matrix_LINE_SEL_Out_c_2), 
            .Matrix_CTRL_Out_c_0(Matrix_CTRL_Out_c_0), .n12311(n12311), 
            .\lastReadRow[4] (lastReadRow[4]), .n10349(n10349), .n12221(n12221), 
            .n13141(n13141), .n87(n87), .\lastReadRow[3] (lastReadRow[3]), 
            .n12342(n12342), .n10350(n10350), .n12284(n12284), .\VRAM_ADDR[6] (VRAM_ADDR[6]), 
            .\VRAM_ADDR[5] (VRAM_ADDR[5]), .\VRAM_ADDR[4] (VRAM_ADDR[4]), 
            .\VRAM_ADDR[3] (VRAM_ADDR[3]), .\VRAM_ADDR[2] (VRAM_ADDR[2]), 
            .\VRAM_ADDR[1] (VRAM_ADDR[1]), .\VRAM_ADDR[0] (VRAM_ADDR[0]), 
            .n3028({n3028}), .n3027({n3027}), .VCC_net(VCC_net), .VRAM_WC(VRAM_WC), 
            .n3035({n3035}), .n3034({n3034}), .n3033({n3033}), .n3032({n3032}), 
            .n3037({n3037}), .n3036({n3036}), .n3030({n3030}), .n3029({n3029}), 
            .n3031({n3031}), .VRAM_DATA({VRAM_DATA}));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(139[6:30])
    LUT4 m1_lut (.Z(n13160)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    
endmodule
//
// Verilog Description of module SRAM
//

module SRAM (lastAddress, LOGIC_CLOCK, lastAddress_31__N_872, n66, SRAM_OE_c, 
            SRAM_WE_c, lastAddress_31__N_785, lastAddress_31__N_845, lastAddress_31__N_857, 
            n55, lastAddress_31__N_786, lastAddress_31__N_781, lastAddress_31__N_777, 
            BUS_DATA_INTERNAL, SRAM_DATA_out_0, SRAM_ADDR_c_0, n12269, 
            lastAddress_31__N_789, lastAddress_31__N_881, n13160, lastAddress_31__N_875, 
            n61, lastAddress_31__N_860, n56, n12057, SRAM_WE_N_704, 
            lastAddress_31__N_782, lastAddress_31__N_827, n33, lastAddress_31__N_836, 
            n48, BUS_DONE_INTERNAL, lastAddress_31__N_787, GND_net, 
            lastAddress_31__N_884, n64, n39, n38, n35, n37, n36, 
            lastAddress_31__N_851, lastAddress_31__N_779, lastAddress_31__N_774, 
            lastAddress_31__N_848, n52, lastAddress_31__N_778, lastAddress_31__N_863, 
            n57, lastAddress_31__N_783, n42, n41, n34, lastAddress_31__N_760, 
            n43, n40, lastAddress_31__N_830, n46, \BUS_ADDR_INTERNAL[18]_derived_1 , 
            lastAddress_31__N_833, n47, n44, n45, lastAddress_31__N_790, 
            lastAddress_31__N_866, n58, n13141, n87, \PWMArray[0][12] , 
            n12221, \MATRIX_data[3] , lastAddress_31__N_784, \PWMArray[0][11] , 
            \MATRIX_data[2] , lastAddress_31__N_839, n49, n12265, n12309, 
            SRAM_DATA_out_1, SRAM_DATA_out_2, SRAM_DATA_out_3, SRAM_DATA_out_4, 
            SRAM_DATA_out_5, SRAM_DATA_out_6, SRAM_DATA_out_7, \BUS_DATA_INTERNAL[8] , 
            SRAM_DATA_out_8, \BUS_DATA_INTERNAL[9] , SRAM_DATA_out_9, 
            \BUS_DATA_INTERNAL[10] , SRAM_DATA_out_10, \BUS_DATA_INTERNAL[11] , 
            SRAM_DATA_out_11, \BUS_DATA_INTERNAL[12] , SRAM_DATA_out_12, 
            \BUS_DATA_INTERNAL[13] , SRAM_DATA_out_13, \BUS_DATA_INTERNAL[14] , 
            SRAM_DATA_out_14, \BUS_DATA_INTERNAL[15] , SRAM_DATA_out_15, 
            SRAM_ADDR_c_1, SRAM_ADDR_c_2, n12253, SRAM_ADDR_c_3, n12264, 
            SRAM_ADDR_c_4, n12259, SRAM_ADDR_c_5, n12247, SRAM_ADDR_c_6, 
            n12252, SRAM_ADDR_c_7, n12263, SRAM_ADDR_c_8, n12250, 
            SRAM_ADDR_c_9, n12271, SRAM_ADDR_c_10, n12268, SRAM_ADDR_c_11, 
            \BUS_addr[11] , SRAM_ADDR_c_12, n12251, SRAM_ADDR_c_13, 
            \BUS_addr[13] , SRAM_ADDR_c_14, \BUS_addr[14] , SRAM_ADDR_c_15, 
            n12270, SRAM_ADDR_c_16, n12262, SRAM_ADDR_c_17, n12329, 
            \PWMArray[0][10] , \MATRIX_data[1] , lastAddress_31__N_788, 
            lastAddress_31__N_878, lastAddress_31__N_869, lastAddress_31__N_780, 
            lastAddress_31__N_854, lastAddress_31__N_776, lastAddress_31__N_842, 
            lastAddress_31__N_775, lastAddress_31__N_773, BUS_DIRECTION_INTERNAL, 
            \BUS_currGrantID[0] , \BUS_currGrantID[1] , n12223, n12217, 
            n12216, n54, MDM_done, n1886, BUS_VALID_N_113, n7, n63, 
            n12227, LOGIC_CLOCK_enable_26, LOGIC_CLOCK_enable_49, n12219, 
            n1184, LOGIC_CLOCK_enable_71, \lastAddress[12] , \lastAddress[10] , 
            n62, n12354, n63_adj_36, PWMArray_0__12__N_110, \lastAddress[16] , 
            n2198, BUS_VALID_N_1118, n12220, n4, \BUS_data[7] , n4_adj_37, 
            \BUS_data[6] , n4_adj_38, \BUS_data[5] , n4_adj_39, \BUS_data[4] , 
            transferMode_3__N_1115, \lastAddress[31] , n12258, \PWMArray[0][9] , 
            \MATRIX_data[0] );
    output [31:0]lastAddress;
    input LOGIC_CLOCK;
    input lastAddress_31__N_872;
    input [31:0]n66;
    output SRAM_OE_c;
    output SRAM_WE_c;
    input lastAddress_31__N_785;
    input lastAddress_31__N_845;
    input lastAddress_31__N_857;
    input n55;
    input lastAddress_31__N_786;
    input lastAddress_31__N_781;
    input lastAddress_31__N_777;
    output [15:0]BUS_DATA_INTERNAL;
    input SRAM_DATA_out_0;
    output SRAM_ADDR_c_0;
    input n12269;
    input lastAddress_31__N_789;
    input lastAddress_31__N_881;
    input n13160;
    input lastAddress_31__N_875;
    input n61;
    input lastAddress_31__N_860;
    input n56;
    input n12057;
    output SRAM_WE_N_704;
    input lastAddress_31__N_782;
    input lastAddress_31__N_827;
    input n33;
    input lastAddress_31__N_836;
    input n48;
    output BUS_DONE_INTERNAL;
    input lastAddress_31__N_787;
    input GND_net;
    input lastAddress_31__N_884;
    input n64;
    input n39;
    input n38;
    input n35;
    input n37;
    input n36;
    input lastAddress_31__N_851;
    input lastAddress_31__N_779;
    input lastAddress_31__N_774;
    input lastAddress_31__N_848;
    input n52;
    input lastAddress_31__N_778;
    input lastAddress_31__N_863;
    input n57;
    input lastAddress_31__N_783;
    input n42;
    input n41;
    input n34;
    input lastAddress_31__N_760;
    input n43;
    input n40;
    input lastAddress_31__N_830;
    input n46;
    input \BUS_ADDR_INTERNAL[18]_derived_1 ;
    input lastAddress_31__N_833;
    input n47;
    input n44;
    input n45;
    input lastAddress_31__N_790;
    input lastAddress_31__N_866;
    input n58;
    input n13141;
    input n87;
    input \PWMArray[0][12] ;
    input n12221;
    output \MATRIX_data[3] ;
    input lastAddress_31__N_784;
    input \PWMArray[0][11] ;
    output \MATRIX_data[2] ;
    input lastAddress_31__N_839;
    input n49;
    input n12265;
    input n12309;
    input SRAM_DATA_out_1;
    input SRAM_DATA_out_2;
    input SRAM_DATA_out_3;
    input SRAM_DATA_out_4;
    input SRAM_DATA_out_5;
    input SRAM_DATA_out_6;
    input SRAM_DATA_out_7;
    output \BUS_DATA_INTERNAL[8] ;
    input SRAM_DATA_out_8;
    output \BUS_DATA_INTERNAL[9] ;
    input SRAM_DATA_out_9;
    output \BUS_DATA_INTERNAL[10] ;
    input SRAM_DATA_out_10;
    output \BUS_DATA_INTERNAL[11] ;
    input SRAM_DATA_out_11;
    output \BUS_DATA_INTERNAL[12] ;
    input SRAM_DATA_out_12;
    output \BUS_DATA_INTERNAL[13] ;
    input SRAM_DATA_out_13;
    output \BUS_DATA_INTERNAL[14] ;
    input SRAM_DATA_out_14;
    output \BUS_DATA_INTERNAL[15] ;
    input SRAM_DATA_out_15;
    output SRAM_ADDR_c_1;
    output SRAM_ADDR_c_2;
    input n12253;
    output SRAM_ADDR_c_3;
    input n12264;
    output SRAM_ADDR_c_4;
    input n12259;
    output SRAM_ADDR_c_5;
    input n12247;
    output SRAM_ADDR_c_6;
    input n12252;
    output SRAM_ADDR_c_7;
    input n12263;
    output SRAM_ADDR_c_8;
    input n12250;
    output SRAM_ADDR_c_9;
    input n12271;
    output SRAM_ADDR_c_10;
    input n12268;
    output SRAM_ADDR_c_11;
    input \BUS_addr[11] ;
    output SRAM_ADDR_c_12;
    input n12251;
    output SRAM_ADDR_c_13;
    input \BUS_addr[13] ;
    output SRAM_ADDR_c_14;
    input \BUS_addr[14] ;
    output SRAM_ADDR_c_15;
    input n12270;
    output SRAM_ADDR_c_16;
    input n12262;
    output SRAM_ADDR_c_17;
    input n12329;
    input \PWMArray[0][10] ;
    output \MATRIX_data[1] ;
    input lastAddress_31__N_788;
    input lastAddress_31__N_878;
    input lastAddress_31__N_869;
    input lastAddress_31__N_780;
    input lastAddress_31__N_854;
    input lastAddress_31__N_776;
    input lastAddress_31__N_842;
    input lastAddress_31__N_775;
    input lastAddress_31__N_773;
    input BUS_DIRECTION_INTERNAL;
    input \BUS_currGrantID[0] ;
    input \BUS_currGrantID[1] ;
    input n12223;
    output n12217;
    output n12216;
    input n54;
    input MDM_done;
    input n1886;
    input BUS_VALID_N_113;
    output n7;
    input n63;
    input n12227;
    input LOGIC_CLOCK_enable_26;
    output LOGIC_CLOCK_enable_49;
    input n12219;
    input n1184;
    output LOGIC_CLOCK_enable_71;
    output \lastAddress[12] ;
    output \lastAddress[10] ;
    input n62;
    input n12354;
    input n63_adj_36;
    output PWMArray_0__12__N_110;
    output \lastAddress[16] ;
    input n2198;
    input BUS_VALID_N_1118;
    output n12220;
    input n4;
    output \BUS_data[7] ;
    input n4_adj_37;
    output \BUS_data[6] ;
    input n4_adj_38;
    output \BUS_data[5] ;
    input n4_adj_39;
    output \BUS_data[4] ;
    output transferMode_3__N_1115;
    output \lastAddress[31] ;
    input n12258;
    input \PWMArray[0][9] ;
    output \MATRIX_data[0] ;
    
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    
    wire n5210, n5209, n5208, LOGIC_CLOCK_enable_2, SRAM_OE_N_961, 
        LOGIC_CLOCK_enable_3, SRAM_WE_N_695, n5213, n5246;
    wire [31:0]n66_c;
    
    wire n5230, n5229, n5266, n5265, n5264, n5245, LOGIC_CLOCK_enable_96, 
        LOGIC_CLOCK_enable_113;
    wire [7:0]state;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(34[8:13])
    wire [7:0]state_7__N_903;
    
    wire n5196, n5206, n5226, n12056, n5225, n5306, n5258, LOGIC_CLOCK_enable_34, 
        n12225, n5205, n10007;
    wire [7:0]n138;
    
    wire n10006, n10005, n10004, n5194, n5291, n5294, n5303, n5297, 
        n5300, n5238, n5237, n5257, n5242, n5241, n5222, n5221, 
        n5282, n5285, n5270, n5269, n5279, n5288, n5262, n5276, 
        n5273, n5193, n5218, n5217, n5261, n5260, n5275, n5268, 
        n5272, n5254, n9692, n9691, n9690;
    wire [15:0]BUS_DATA_INTERNAL_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(30[8:25])
    wire [7:0]state_7__N_911;
    
    wire n5200, n5204, n5212, n5216, n5220, n5224, n5228, n5232, 
        n5236, n5240, n5244, n5248, n5252, n5256, n5278, n5281, 
        n5284, n5287, n5290, n5293, n5296, n5299, n5302, n5305, 
        n5253, n5234, n9689, n9688, n9687;
    wire [31:0]lastAddress_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(29[8:19])
    
    wire n5198, n5197, n5202, n12110, n12310, n12111, n12257, 
        n12353, n12283, n5214, n5233, n5192, n5201, n5250, n5249, 
        n9686, n12282, n10, n12341;
    
    LUT4 i2614_3_lut (.A(n5210), .B(n5209), .C(n5208), .Z(lastAddress[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2614_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i4_2612_2613_reset (.D(n66[4]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_872), .Q(n5210)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i4_2612_2613_reset.GSR = "DISABLED";
    FD1P3AY SRAM_OE_INT_225 (.D(SRAM_OE_N_961), .SP(LOGIC_CLOCK_enable_2), 
            .CK(LOGIC_CLOCK), .Q(SRAM_OE_c)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_OE_INT_225.GSR = "ENABLED";
    FD1P3AY SRAM_WE_INT_224 (.D(SRAM_WE_N_695), .SP(LOGIC_CLOCK_enable_3), 
            .CK(LOGIC_CLOCK), .Q(SRAM_WE_c)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_WE_INT_224.GSR = "ENABLED";
    FD1S3BX lastAddress_i0_i5_2616_2617_set (.D(n66[5]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_785), .Q(n5213)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i5_2616_2617_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i13_2648_2649_reset (.D(n66_c[13]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_845), .Q(n5246)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i13_2648_2649_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i9_2632_2633_reset (.D(n55), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_857), .Q(n5230)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i9_2632_2633_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i4_2612_2613_set (.D(n66[4]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_786), .Q(n5209)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i4_2612_2613_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i9_2632_2633_set (.D(n55), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_781), .Q(n5229)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i9_2632_2633_set.GSR = "DISABLED";
    LUT4 i2670_3_lut (.A(n5266), .B(n5265), .C(n5264), .Z(lastAddress[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2670_3_lut.init = 16'hcaca;
    FD1S3BX lastAddress_i0_i13_2648_2649_set (.D(n66_c[13]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_777), .Q(n5245)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i13_2648_2649_set.GSR = "DISABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i0 (.D(SRAM_DATA_out_0), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i0.GSR = "ENABLED";
    FD1P3AX SRAM_ADDR_i0_i1 (.D(n12269), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i1.GSR = "DISABLED";
    FD1S3AX state_i0 (.D(state_7__N_903[0]), .CK(LOGIC_CLOCK), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i0.GSR = "ENABLED";
    FD1S1D i2599 (.D(n13160), .CK(lastAddress_31__N_789), .CD(lastAddress_31__N_881), 
           .Q(n5196));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2599.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i3_2608_2609_reset (.D(n61), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_875), .Q(n5206)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i3_2608_2609_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i8_2628_2629_reset (.D(n56), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_860), .Q(n5226)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i8_2628_2629_reset.GSR = "DISABLED";
    PFUMX i8968 (.BLUT(n12057), .ALUT(n12056), .C0(SRAM_WE_N_704), .Z(state_7__N_903[0]));
    FD1S3BX lastAddress_i0_i8_2628_2629_set (.D(n56), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_782), .Q(n5225)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i8_2628_2629_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i31_2708_2709_reset (.D(n33), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5306)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i31_2708_2709_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i16_2660_2661_reset (.D(n48), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_836), .Q(n5258)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i16_2660_2661_reset.GSR = "DISABLED";
    FD1P3IX BUS_DONE_INTERNAL_123 (.D(n13160), .SP(LOGIC_CLOCK_enable_34), 
            .CD(n12225), .CK(LOGIC_CLOCK), .Q(BUS_DONE_INTERNAL)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DONE_INTERNAL_123.GSR = "ENABLED";
    FD1S3BX lastAddress_i0_i3_2608_2609_set (.D(n61), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_787), .Q(n5205)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i3_2608_2609_set.GSR = "DISABLED";
    CCU2D add_90_9 (.A0(state[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10007), 
          .S0(n138[7]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_90_9.INIT0 = 16'h5aaa;
    defparam add_90_9.INIT1 = 16'h0000;
    defparam add_90_9.INJECT1_0 = "NO";
    defparam add_90_9.INJECT1_1 = "NO";
    CCU2D add_90_7 (.A0(state[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(state[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10006), 
          .COUT(n10007), .S0(n138[5]), .S1(n138[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_90_7.INIT0 = 16'h5aaa;
    defparam add_90_7.INIT1 = 16'h5aaa;
    defparam add_90_7.INJECT1_0 = "NO";
    defparam add_90_7.INJECT1_1 = "NO";
    CCU2D add_90_5 (.A0(state[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(state[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10005), 
          .COUT(n10006), .S0(n138[3]), .S1(n138[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_90_5.INIT0 = 16'h5aaa;
    defparam add_90_5.INIT1 = 16'h5aaa;
    defparam add_90_5.INJECT1_0 = "NO";
    defparam add_90_5.INJECT1_1 = "NO";
    CCU2D add_90_3 (.A0(state[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(state[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10004), 
          .COUT(n10005), .S0(n138[1]), .S1(n138[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_90_3.INIT0 = 16'h5aaa;
    defparam add_90_3.INIT1 = 16'h5aaa;
    defparam add_90_3.INJECT1_0 = "NO";
    defparam add_90_3.INJECT1_1 = "NO";
    FD1S3DX lastAddress_i0_i0_2596_2597_reset (.D(n64), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_884), .Q(n5194)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i0_2596_2597_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i25_2693_2694_reset (.D(n39), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5291)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i25_2693_2694_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i26_2696_2697_reset (.D(n38), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5294)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i26_2696_2697_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i29_2705_2706_reset (.D(n35), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5303)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i29_2705_2706_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i27_2699_2700_reset (.D(n37), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5297)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i27_2699_2700_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i28_2702_2703_reset (.D(n36), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5300)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i28_2702_2703_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i11_2640_2641_reset (.D(n66_c[11]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_851), .Q(n5238)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i11_2640_2641_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i11_2640_2641_set (.D(n66_c[11]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_779), .Q(n5237)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i11_2640_2641_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i16_2660_2661_set (.D(n48), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_774), .Q(n5257)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i16_2660_2661_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i12_2644_2645_reset (.D(n52), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_848), .Q(n5242)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i12_2644_2645_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i12_2644_2645_set (.D(n52), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_778), .Q(n5241)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i12_2644_2645_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i7_2624_2625_reset (.D(n57), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_863), .Q(n5222)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i7_2624_2625_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i7_2624_2625_set (.D(n57), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_783), .Q(n5221)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i7_2624_2625_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i22_2684_2685_reset (.D(n42), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5282)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i22_2684_2685_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i23_2687_2688_reset (.D(n41), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5285)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i23_2687_2688_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i30_2672_2673_reset (.D(n34), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5270)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i30_2672_2673_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i30_2672_2673_set (.D(n34), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5269)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i30_2672_2673_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i21_2681_2682_reset (.D(n43), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5279)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i21_2681_2682_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i24_2690_2691_reset (.D(n40), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5288)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i24_2690_2691_reset.GSR = "DISABLED";
    CCU2D add_90_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(state[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n10004), 
          .S1(n138[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_90_1.INIT0 = 16'hF000;
    defparam add_90_1.INIT1 = 16'h5555;
    defparam add_90_1.INJECT1_0 = "NO";
    defparam add_90_1.INJECT1_1 = "NO";
    FD1S3DX lastAddress_i0_i18_2668_2669_reset (.D(n46), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_830), .Q(n5266)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i18_2668_2669_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i18_2668_2669_set (.D(n46), .CK(LOGIC_CLOCK), 
            .PD(\BUS_ADDR_INTERNAL[18]_derived_1 ), .Q(n5265)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i18_2668_2669_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i17_2664_2665_reset (.D(n47), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_833), .Q(n5262)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i17_2664_2665_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i20_2678_2679_reset (.D(n44), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5276)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i20_2678_2679_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i19_2675_2676_reset (.D(n45), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_827), .Q(n5273)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i19_2675_2676_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i0_2596_2597_set (.D(n64), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_790), .Q(n5193)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i0_2596_2597_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i6_2620_2621_reset (.D(n58), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_866), .Q(n5218)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i6_2620_2621_reset.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n13141), .B(n87), .C(\PWMArray[0][12] ), 
         .D(n12221), .Z(\MATRIX_data[3] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    FD1S3BX lastAddress_i0_i6_2620_2621_set (.D(n58), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_784), .Q(n5217)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i6_2620_2621_set.GSR = "DISABLED";
    LUT4 i2666_3_lut (.A(n5262), .B(n5261), .C(n5260), .Z(lastAddress[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2666_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_182 (.A(n13141), .B(n87), .C(\PWMArray[0][11] ), 
         .D(n12221), .Z(\MATRIX_data[2] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_182.init = 16'h1000;
    LUT4 i2680_3_lut (.A(n5276), .B(n5275), .C(n5268), .Z(lastAddress[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2680_3_lut.init = 16'hcaca;
    LUT4 i2677_3_lut (.A(n5273), .B(n5272), .C(n5268), .Z(lastAddress[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2677_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i15_2656_2657_reset (.D(n49), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_839), .Q(n5254)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i15_2656_2657_reset.GSR = "DISABLED";
    CCU2D lastAddress_31__I_0_299_32 (.A0(lastAddress[22]), .B0(lastAddress[21]), 
          .C0(lastAddress[20]), .D0(lastAddress[19]), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n9692), .S1(SRAM_WE_N_704));
    defparam lastAddress_31__I_0_299_32.INIT0 = 16'h8001;
    defparam lastAddress_31__I_0_299_32.INIT1 = 16'hFFFF;
    defparam lastAddress_31__I_0_299_32.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_32.INJECT1_1 = "NO";
    CCU2D lastAddress_31__I_0_299_31 (.A0(lastAddress[28]), .B0(lastAddress[27]), 
          .C0(lastAddress[26]), .D0(lastAddress[25]), .A1(lastAddress[25]), 
          .B1(lastAddress[24]), .C1(lastAddress[23]), .D1(lastAddress[22]), 
          .CIN(n9691), .COUT(n9692));
    defparam lastAddress_31__I_0_299_31.INIT0 = 16'h8001;
    defparam lastAddress_31__I_0_299_31.INIT1 = 16'h8001;
    defparam lastAddress_31__I_0_299_31.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_31.INJECT1_1 = "YES";
    CCU2D lastAddress_31__I_0_299_29 (.A0(n12265), .B0(lastAddress[1]), 
          .C0(n12269), .D0(lastAddress[0]), .A1(n12309), .B1(lastAddress[30]), 
          .C1(lastAddress[29]), .D1(lastAddress[28]), .CIN(n9690), .COUT(n9691));
    defparam lastAddress_31__I_0_299_29.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_299_29.INIT1 = 16'h8001;
    defparam lastAddress_31__I_0_299_29.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_29.INJECT1_1 = "YES";
    FD1P3AX BUS_DATA_INTERNAL_i0_i1 (.D(SRAM_DATA_out_1), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i1.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i2 (.D(SRAM_DATA_out_2), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i2.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i3 (.D(SRAM_DATA_out_3), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i3.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i4 (.D(SRAM_DATA_out_4), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL_c[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i4.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i5 (.D(SRAM_DATA_out_5), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL_c[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i5.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i6 (.D(SRAM_DATA_out_6), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL_c[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i6.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i7 (.D(SRAM_DATA_out_7), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(BUS_DATA_INTERNAL_c[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i7.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i8 (.D(SRAM_DATA_out_8), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i8.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i9 (.D(SRAM_DATA_out_9), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i9.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i10 (.D(SRAM_DATA_out_10), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i10.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i11 (.D(SRAM_DATA_out_11), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i11.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i12 (.D(SRAM_DATA_out_12), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i12.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i13 (.D(SRAM_DATA_out_13), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[13] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i13.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i14 (.D(SRAM_DATA_out_14), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[14] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i14.GSR = "ENABLED";
    FD1P3AX BUS_DATA_INTERNAL_i0_i15 (.D(SRAM_DATA_out_15), .SP(LOGIC_CLOCK_enable_96), 
            .CK(LOGIC_CLOCK), .Q(\BUS_DATA_INTERNAL[15] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam BUS_DATA_INTERNAL_i0_i15.GSR = "ENABLED";
    FD1P3AX SRAM_ADDR_i0_i2 (.D(n12265), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i2.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i3 (.D(n12253), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i3.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i4 (.D(n12264), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i4.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i5 (.D(n12259), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i5.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i6 (.D(n12247), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i6.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i7 (.D(n12252), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i7.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i8 (.D(n12263), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i8.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i9 (.D(n12250), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i9.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i10 (.D(n12271), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_9)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i10.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i11 (.D(n12268), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_10)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i11.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i12 (.D(\BUS_addr[11] ), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(SRAM_ADDR_c_11)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i12.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i13 (.D(n12251), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_12)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i13.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i14 (.D(\BUS_addr[13] ), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(SRAM_ADDR_c_13)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i14.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i15 (.D(\BUS_addr[14] ), .SP(LOGIC_CLOCK_enable_113), 
            .CK(LOGIC_CLOCK), .Q(SRAM_ADDR_c_14)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i15.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i16 (.D(n12270), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_15)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i16.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i17 (.D(n12262), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_16)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i17.GSR = "DISABLED";
    FD1P3AX SRAM_ADDR_i0_i18 (.D(n12329), .SP(LOGIC_CLOCK_enable_113), .CK(LOGIC_CLOCK), 
            .Q(SRAM_ADDR_c_17)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam SRAM_ADDR_i0_i18.GSR = "DISABLED";
    FD1S3AX state_i1 (.D(state_7__N_903[1]), .CK(LOGIC_CLOCK), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_183 (.A(n13141), .B(n87), .C(\PWMArray[0][10] ), 
         .D(n12221), .Z(\MATRIX_data[1] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_183.init = 16'h1000;
    FD1S3AX state_i2 (.D(state_7__N_903[2]), .CK(LOGIC_CLOCK), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i3 (.D(state_7__N_903[3]), .CK(LOGIC_CLOCK), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i3.GSR = "ENABLED";
    FD1S3AX state_i4 (.D(state_7__N_903[4]), .CK(LOGIC_CLOCK), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i4.GSR = "ENABLED";
    FD1S3IX state_i5 (.D(state_7__N_911[5]), .CK(LOGIC_CLOCK), .CD(n12225), 
            .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i5.GSR = "ENABLED";
    FD1S3IX state_i6 (.D(state_7__N_911[6]), .CK(LOGIC_CLOCK), .CD(n12225), 
            .Q(state[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i6.GSR = "ENABLED";
    FD1S3IX state_i7 (.D(state_7__N_911[7]), .CK(LOGIC_CLOCK), .CD(n12225), 
            .Q(state[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam state_i7.GSR = "ENABLED";
    FD1S1D i2603 (.D(n13160), .CK(lastAddress_31__N_788), .CD(lastAddress_31__N_878), 
           .Q(n5200));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2603.GSR = "DISABLED";
    FD1S1D i2607 (.D(n13160), .CK(lastAddress_31__N_787), .CD(lastAddress_31__N_875), 
           .Q(n5204));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2607.GSR = "DISABLED";
    FD1S1D i2611 (.D(n13160), .CK(lastAddress_31__N_786), .CD(lastAddress_31__N_872), 
           .Q(n5208));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2611.GSR = "DISABLED";
    FD1S1D i2615 (.D(n13160), .CK(lastAddress_31__N_785), .CD(lastAddress_31__N_869), 
           .Q(n5212));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2615.GSR = "DISABLED";
    FD1S1D i2619 (.D(n13160), .CK(lastAddress_31__N_784), .CD(lastAddress_31__N_866), 
           .Q(n5216));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2619.GSR = "DISABLED";
    FD1S1D i2623 (.D(n13160), .CK(lastAddress_31__N_783), .CD(lastAddress_31__N_863), 
           .Q(n5220));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2623.GSR = "DISABLED";
    FD1S1D i2627 (.D(n13160), .CK(lastAddress_31__N_782), .CD(lastAddress_31__N_860), 
           .Q(n5224));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2627.GSR = "DISABLED";
    FD1S1D i2631 (.D(n13160), .CK(lastAddress_31__N_781), .CD(lastAddress_31__N_857), 
           .Q(n5228));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2631.GSR = "DISABLED";
    FD1S1D i2635 (.D(n13160), .CK(lastAddress_31__N_780), .CD(lastAddress_31__N_854), 
           .Q(n5232));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2635.GSR = "DISABLED";
    FD1S1D i2639 (.D(n13160), .CK(lastAddress_31__N_779), .CD(lastAddress_31__N_851), 
           .Q(n5236));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2639.GSR = "DISABLED";
    FD1S1D i2643 (.D(n13160), .CK(lastAddress_31__N_778), .CD(lastAddress_31__N_848), 
           .Q(n5240));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2643.GSR = "DISABLED";
    FD1S1D i2647 (.D(n13160), .CK(lastAddress_31__N_777), .CD(lastAddress_31__N_845), 
           .Q(n5244));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2647.GSR = "DISABLED";
    FD1S1D i2651 (.D(n13160), .CK(lastAddress_31__N_776), .CD(lastAddress_31__N_842), 
           .Q(n5248));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2651.GSR = "DISABLED";
    FD1S1D i2655 (.D(n13160), .CK(lastAddress_31__N_775), .CD(lastAddress_31__N_839), 
           .Q(n5252));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2655.GSR = "DISABLED";
    FD1S1D i2659 (.D(n13160), .CK(lastAddress_31__N_774), .CD(lastAddress_31__N_836), 
           .Q(n5256));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2659.GSR = "DISABLED";
    FD1S1D i2663 (.D(n13160), .CK(lastAddress_31__N_773), .CD(lastAddress_31__N_833), 
           .Q(n5260));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2663.GSR = "DISABLED";
    FD1S1D i2667 (.D(n13160), .CK(\BUS_ADDR_INTERNAL[18]_derived_1 ), .CD(lastAddress_31__N_830), 
           .Q(n5264));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2667.GSR = "DISABLED";
    FD1S1D i2671 (.D(n13160), .CK(lastAddress_31__N_760), .CD(lastAddress_31__N_827), 
           .Q(n5268));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2671.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i20_2678_2679_set (.D(n44), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5275)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i20_2678_2679_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i21_2681_2682_set (.D(n43), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5278)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i21_2681_2682_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i22_2684_2685_set (.D(n42), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5281)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i22_2684_2685_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i23_2687_2688_set (.D(n41), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5284)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i23_2687_2688_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i24_2690_2691_set (.D(n40), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5287)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i24_2690_2691_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i25_2693_2694_set (.D(n39), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5290)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i25_2693_2694_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i26_2696_2697_set (.D(n38), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5293)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i26_2696_2697_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i27_2699_2700_set (.D(n37), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5296)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i27_2699_2700_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i28_2702_2703_set (.D(n36), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5299)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i28_2702_2703_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i29_2705_2706_set (.D(n35), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5302)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i29_2705_2706_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i31_2708_2709_set (.D(n33), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5305)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i31_2708_2709_set.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i19_2675_2676_set (.D(n45), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_760), .Q(n5272)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i19_2675_2676_set.GSR = "DISABLED";
    LUT4 OUT_ENABLE_I_0_3_lut_rep_191_4_lut_4_lut_3_lut_4_lut_4_lut (.A(BUS_DIRECTION_INTERNAL), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .D(n12223), 
         .Z(n12217)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam OUT_ENABLE_I_0_3_lut_rep_191_4_lut_4_lut_3_lut_4_lut_4_lut.init = 16'h3c10;
    LUT4 i1603_2_lut_rep_190_4_lut_4_lut_4_lut_4_lut_4_lut (.A(BUS_DIRECTION_INTERNAL), 
         .B(\BUS_currGrantID[0] ), .C(\BUS_currGrantID[1] ), .Z(n12216)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1603_2_lut_rep_190_4_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h1010;
    LUT4 i2658_3_lut (.A(n5254), .B(n5253), .C(n5252), .Z(lastAddress[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2658_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i10_2636_2637_reset (.D(n54), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_854), .Q(n5234)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i10_2636_2637_reset.GSR = "DISABLED";
    CCU2D lastAddress_31__I_0_299_27 (.A0(n12247), .B0(lastAddress[5]), 
          .C0(n12259), .D0(lastAddress[4]), .A1(n12264), .B1(lastAddress[3]), 
          .C1(n12253), .D1(lastAddress[2]), .CIN(n9689), .COUT(n9690));
    defparam lastAddress_31__I_0_299_27.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_299_27.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_299_27.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_27.INJECT1_1 = "YES";
    CCU2D lastAddress_31__I_0_299_25 (.A0(n12271), .B0(lastAddress[9]), 
          .C0(n12250), .D0(lastAddress[8]), .A1(n12263), .B1(lastAddress[7]), 
          .C1(n12252), .D1(lastAddress[6]), .CIN(n9688), .COUT(n9689));
    defparam lastAddress_31__I_0_299_25.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_299_25.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_299_25.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_25.INJECT1_1 = "YES";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_184 (.A(n13141), .B(MDM_done), .C(n1886), 
         .D(BUS_VALID_N_113), .Z(n7)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_184.init = 16'hcdcc;
    FD1S3BX lastAddress_i0_i15_2656_2657_set (.D(n49), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_775), .Q(n5253)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i15_2656_2657_set.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_4_lut (.A(n13141), .B(n63), .C(n12227), .D(LOGIC_CLOCK_enable_26), 
         .Z(LOGIC_CLOCK_enable_49)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n13141), .B(n12219), .C(n1184), 
         .D(LOGIC_CLOCK_enable_26), .Z(LOGIC_CLOCK_enable_71)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h0002;
    CCU2D lastAddress_31__I_0_299_23 (.A0(\BUS_addr[13] ), .B0(lastAddress_c[13]), 
          .C0(n12251), .D0(\lastAddress[12] ), .A1(\BUS_addr[11] ), .B1(lastAddress_c[11]), 
          .C1(n12268), .D1(\lastAddress[10] ), .CIN(n9687), .COUT(n9688));
    defparam lastAddress_31__I_0_299_23.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_299_23.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_299_23.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_23.INJECT1_1 = "YES";
    LUT4 i2602_3_lut (.A(n5198), .B(n5197), .C(n5196), .Z(lastAddress[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2602_3_lut.init = 16'hcaca;
    FD1S3DX lastAddress_i0_i2_2604_2605_reset (.D(n62), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_878), .Q(n5202)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i2_2604_2605_reset.GSR = "DISABLED";
    LUT4 state_7__N_919_0__bdd_3_lut (.A(n13141), .B(state[4]), .C(state[5]), 
         .Z(n12110)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam state_7__N_919_0__bdd_3_lut.init = 16'hfefe;
    LUT4 n12110_bdd_3_lut (.A(n12110), .B(n138[4]), .C(n12310), .Z(n12111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n12110_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_231_3_lut (.A(n12310), .B(state[4]), .C(state[5]), 
         .Z(n12257)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(94[10:23])
    defparam i1_2_lut_rep_231_3_lut.init = 16'hfefe;
    PFUMX i9057 (.BLUT(n12353), .ALUT(n12354), .C0(n12310), .Z(LOGIC_CLOCK_enable_3));
    LUT4 i8599_2_lut_3_lut_3_lut_4_lut_3_lut_4_lut (.A(n12310), .B(state[4]), 
         .C(SRAM_WE_N_704), .D(state[5]), .Z(SRAM_WE_N_695)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(94[10:23])
    defparam i8599_2_lut_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_rep_257 (.A(n12310), .B(state[4]), .C(state[5]), .Z(n12283)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(78[10:23])
    defparam i2_3_lut_rep_257.init = 16'hfbfb;
    LUT4 i8603_3_lut_4_lut_4_lut (.A(n13141), .B(n12283), .C(SRAM_WE_N_704), 
         .D(n12257), .Z(LOGIC_CLOCK_enable_2)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i8603_3_lut_4_lut_4_lut.init = 16'h3555;
    FD1S3DX lastAddress_i0_i5_2616_2617_reset (.D(n66[5]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_869), .Q(n5214)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i5_2616_2617_reset.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i10_2636_2637_set (.D(n54), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_780), .Q(n5233)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i10_2636_2637_set.GSR = "DISABLED";
    FD1S1D i2595 (.D(n13160), .CK(lastAddress_31__N_790), .CD(lastAddress_31__N_884), 
           .Q(n5192));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2595.GSR = "DISABLED";
    FD1S3BX lastAddress_i0_i2_2604_2605_set (.D(n62), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_788), .Q(n5201)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i2_2604_2605_set.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i14_2652_2653_reset (.D(n66_c[14]), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_842), .Q(n5250)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i14_2652_2653_reset.GSR = "DISABLED";
    FD1S3DX lastAddress_i0_i1_2600_2601_reset (.D(n63_adj_36), .CK(LOGIC_CLOCK), 
            .CD(lastAddress_31__N_881), .Q(n5198)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i1_2600_2601_reset.GSR = "DISABLED";
    LUT4 i2638_3_lut (.A(n5234), .B(n5233), .C(n5232), .Z(\lastAddress[10] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2638_3_lut.init = 16'hcaca;
    LUT4 i2606_3_lut (.A(n5202), .B(n5201), .C(n5200), .Z(lastAddress[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2606_3_lut.init = 16'hcaca;
    LUT4 PWMArray_0__12__I_6_2_lut_3_lut_3_lut (.A(n13141), .B(n1886), .C(BUS_VALID_N_113), 
         .Z(PWMArray_0__12__N_110)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam PWMArray_0__12__I_6_2_lut_3_lut_3_lut.init = 16'hdfdf;
    FD1S3BX lastAddress_i0_i14_2652_2653_set (.D(n66_c[14]), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_776), .Q(n5249)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i14_2652_2653_set.GSR = "DISABLED";
    LUT4 i2622_3_lut (.A(n5218), .B(n5217), .C(n5216), .Z(lastAddress[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2622_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n12257), .B(SRAM_WE_N_704), .C(n12310), .D(n138[1]), 
         .Z(state_7__N_903[1])) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf777;
    LUT4 i1_3_lut_4_lut_adj_185 (.A(n12257), .B(SRAM_WE_N_704), .C(n12310), 
         .D(n138[2]), .Z(state_7__N_903[2])) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_185.init = 16'hf777;
    LUT4 i2654_3_lut (.A(n5250), .B(n5249), .C(n5248), .Z(lastAddress_c[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2654_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_186 (.A(n12257), .B(SRAM_WE_N_704), .C(n12310), 
         .D(n138[3]), .Z(state_7__N_903[3])) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_186.init = 16'hf777;
    CCU2D lastAddress_31__I_0_299_21 (.A0(n12329), .B0(lastAddress[17]), 
          .C0(n12262), .D0(\lastAddress[16] ), .A1(n12270), .B1(lastAddress[15]), 
          .C1(\BUS_addr[14] ), .D1(lastAddress_c[14]), .CIN(n9686), .COUT(n9687));
    defparam lastAddress_31__I_0_299_21.INIT0 = 16'h9009;
    defparam lastAddress_31__I_0_299_21.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_299_21.INJECT1_0 = "YES";
    defparam lastAddress_31__I_0_299_21.INJECT1_1 = "YES";
    LUT4 SRAM_WE_I_89_1_lut_rep_199 (.A(SRAM_WE_N_704), .Z(n12225)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[7:38])
    defparam SRAM_WE_I_89_1_lut_rep_199.init = 16'h5555;
    LUT4 i2610_3_lut (.A(n5206), .B(n5205), .C(n5204), .Z(lastAddress[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2610_3_lut.init = 16'hcaca;
    LUT4 i2630_3_lut (.A(n5226), .B(n5225), .C(n5224), .Z(lastAddress[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2630_3_lut.init = 16'hcaca;
    LUT4 BUS_VALID_I_0_2_lut_rep_194_3_lut_3_lut (.A(n13141), .B(n2198), 
         .C(BUS_VALID_N_1118), .Z(n12220)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam BUS_VALID_I_0_2_lut_rep_194_3_lut_3_lut.init = 16'h1010;
    LUT4 lastAddress_i1_i12_3_lut_3_lut (.A(SRAM_WE_N_704), .B(\BUS_addr[11] ), 
         .C(lastAddress_c[11]), .Z(n66_c[11])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[7:38])
    defparam lastAddress_i1_i12_3_lut_3_lut.init = 16'he4e4;
    LUT4 i2634_3_lut (.A(n5230), .B(n5229), .C(n5228), .Z(lastAddress[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2634_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_4_lut_adj_187 (.A(n13141), .B(BUS_DATA_INTERNAL_c[7]), 
         .C(n4), .D(\BUS_ADDR_INTERNAL[18]_derived_1 ), .Z(\BUS_data[7] )) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i2_3_lut_4_lut_4_lut_adj_187.init = 16'hf0f4;
    LUT4 i2_3_lut_4_lut_4_lut_adj_188 (.A(n13141), .B(BUS_DATA_INTERNAL_c[6]), 
         .C(n4_adj_37), .D(\BUS_ADDR_INTERNAL[18]_derived_1 ), .Z(\BUS_data[6] )) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i2_3_lut_4_lut_4_lut_adj_188.init = 16'hf0f4;
    LUT4 i2_3_lut_4_lut_4_lut_adj_189 (.A(n13141), .B(BUS_DATA_INTERNAL_c[5]), 
         .C(n4_adj_38), .D(\BUS_ADDR_INTERNAL[18]_derived_1 ), .Z(\BUS_data[5] )) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i2_3_lut_4_lut_4_lut_adj_189.init = 16'hf0f4;
    LUT4 i2_3_lut_4_lut_4_lut_adj_190 (.A(n13141), .B(BUS_DATA_INTERNAL_c[4]), 
         .C(n4_adj_39), .D(\BUS_ADDR_INTERNAL[18]_derived_1 ), .Z(\BUS_data[4] )) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i2_3_lut_4_lut_4_lut_adj_190.init = 16'hf0f4;
    LUT4 transferMode_3__I_108_2_lut_3_lut_3_lut (.A(n13141), .B(n2198), 
         .C(BUS_VALID_N_1118), .Z(transferMode_3__N_1115)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam transferMode_3__I_108_2_lut_3_lut_3_lut.init = 16'hdfdf;
    LUT4 i2710_3_lut (.A(n5306), .B(n5305), .C(n5268), .Z(\lastAddress[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2710_3_lut.init = 16'hcaca;
    LUT4 i4983_3_lut_4_lut_4_lut_else_2_lut (.A(n13141), .B(SRAM_WE_N_704), 
         .C(state[4]), .D(state[5]), .Z(n12353)) /* synthesis lut_function=(!(A (B (C))+!A ((C+!(D))+!B))) */ ;
    defparam i4983_3_lut_4_lut_4_lut_else_2_lut.init = 16'h2e2a;
    LUT4 lastAddress_i1_i15_3_lut_3_lut (.A(SRAM_WE_N_704), .B(\BUS_addr[14] ), 
         .C(lastAddress_c[14]), .Z(n66_c[14])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[7:38])
    defparam lastAddress_i1_i15_3_lut_3_lut.init = 16'he4e4;
    FD1S3BX lastAddress_i0_i1_2600_2601_set (.D(n63_adj_36), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_789), .Q(n5197)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i1_2600_2601_set.GSR = "DISABLED";
    LUT4 lastAddress_i1_i14_3_lut (.A(lastAddress_c[13]), .B(\BUS_addr[13] ), 
         .C(SRAM_WE_N_704), .Z(n66_c[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i1_i14_3_lut.init = 16'hacac;
    FD1S3BX lastAddress_i0_i17_2664_2665_set (.D(n47), .CK(LOGIC_CLOCK), 
            .PD(lastAddress_31__N_773), .Q(n5261)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=23, LSE_LLINE=192, LSE_RLINE=192 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam lastAddress_i0_i17_2664_2665_set.GSR = "DISABLED";
    LUT4 i2662_3_lut (.A(n5258), .B(n5257), .C(n5256), .Z(\lastAddress[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2662_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(state[5]), .B(n12282), .C(n12283), .D(SRAM_WE_N_704), 
         .Z(LOGIC_CLOCK_enable_96)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0e00;
    LUT4 i8684_2_lut_2_lut_3_lut_4_lut (.A(state[5]), .B(n12282), .C(n12258), 
         .D(SRAM_WE_N_704), .Z(LOGIC_CLOCK_enable_113)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i8684_2_lut_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i8722_2_lut_3_lut_4_lut_4_lut (.A(n12283), .B(SRAM_WE_N_704), .C(n12282), 
         .D(state[5]), .Z(SRAM_OE_N_961)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i8722_2_lut_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 i5_3_lut_rep_284 (.A(state[1]), .B(n10), .C(state[2]), .Z(n12310)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut_rep_284.init = 16'hfefe;
    LUT4 i4_4_lut (.A(state[0]), .B(state[3]), .C(state[6]), .D(state[7]), 
         .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_256_4_lut (.A(state[1]), .B(n10), .C(state[2]), 
         .D(state[4]), .Z(n12282)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_256_4_lut.init = 16'hfffe;
    LUT4 i8688_2_lut_2_lut_4_lut (.A(state[1]), .B(n10), .C(state[2]), 
         .D(n12341), .Z(LOGIC_CLOCK_enable_34)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i8688_2_lut_2_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_4_lut (.A(state[1]), .B(n10), .C(state[2]), .D(n138[6]), 
         .Z(state_7__N_911[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_4_lut_adj_191 (.A(state[1]), .B(n10), .C(state[2]), 
         .D(n138[7]), .Z(state_7__N_911[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_191.init = 16'hfe00;
    LUT4 i2618_3_lut (.A(n5214), .B(n5213), .C(n5212), .Z(lastAddress[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2618_3_lut.init = 16'hcaca;
    LUT4 i2598_3_lut (.A(n5194), .B(n5193), .C(n5192), .Z(lastAddress[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2598_3_lut.init = 16'hcaca;
    CCU2D lastAddress_31__I_0_299_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n12309), .B1(\lastAddress[31] ), .C1(\BUS_ADDR_INTERNAL[18]_derived_1 ), 
          .D1(lastAddress[18]), .COUT(n9686));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(66[12:37])
    defparam lastAddress_31__I_0_299_0.INIT0 = 16'hF000;
    defparam lastAddress_31__I_0_299_0.INIT1 = 16'h9009;
    defparam lastAddress_31__I_0_299_0.INJECT1_0 = "NO";
    defparam lastAddress_31__I_0_299_0.INJECT1_1 = "YES";
    LUT4 i2695_3_lut (.A(n5291), .B(n5290), .C(n5268), .Z(lastAddress[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2695_3_lut.init = 16'hcaca;
    LUT4 i2698_3_lut (.A(n5294), .B(n5293), .C(n5268), .Z(lastAddress[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2698_3_lut.init = 16'hcaca;
    LUT4 i2707_3_lut (.A(n5303), .B(n5302), .C(n5268), .Z(lastAddress[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2707_3_lut.init = 16'hcaca;
    LUT4 i2701_3_lut (.A(n5297), .B(n5296), .C(n5268), .Z(lastAddress[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2701_3_lut.init = 16'hcaca;
    LUT4 i2704_3_lut (.A(n5300), .B(n5299), .C(n5268), .Z(lastAddress[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2704_3_lut.init = 16'hcaca;
    LUT4 i2642_3_lut (.A(n5238), .B(n5237), .C(n5236), .Z(lastAddress_c[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2642_3_lut.init = 16'hcaca;
    LUT4 state_7__N_919_0__bdd_4_lut (.A(n13141), .B(n12257), .C(n12310), 
         .D(n138[0]), .Z(n12056)) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;
    defparam state_7__N_919_0__bdd_4_lut.init = 16'hf111;
    LUT4 i2646_3_lut (.A(n5242), .B(n5241), .C(n5240), .Z(\lastAddress[12] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2646_3_lut.init = 16'hcaca;
    LUT4 i2626_3_lut (.A(n5222), .B(n5221), .C(n5220), .Z(lastAddress[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2626_3_lut.init = 16'hcaca;
    LUT4 i2686_3_lut (.A(n5282), .B(n5281), .C(n5268), .Z(lastAddress[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2686_3_lut.init = 16'hcaca;
    LUT4 i2689_3_lut (.A(n5285), .B(n5284), .C(n5268), .Z(lastAddress[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2689_3_lut.init = 16'hcaca;
    LUT4 i2674_3_lut (.A(n5270), .B(n5269), .C(n5268), .Z(lastAddress[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2674_3_lut.init = 16'hcaca;
    LUT4 i2683_3_lut (.A(n5279), .B(n5278), .C(n5268), .Z(lastAddress[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2683_3_lut.init = 16'hcaca;
    PFUMX i8992 (.BLUT(n13141), .ALUT(n12111), .C0(SRAM_WE_N_704), .Z(state_7__N_903[4]));
    LUT4 i2692_3_lut (.A(n5288), .B(n5287), .C(n5268), .Z(lastAddress[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2692_3_lut.init = 16'hcaca;
    LUT4 i8114_2_lut_rep_315 (.A(state[4]), .B(state[5]), .Z(n12341)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8114_2_lut_rep_315.init = 16'heeee;
    LUT4 i14_3_lut_4_lut (.A(state[4]), .B(state[5]), .C(n12310), .D(n138[5]), 
         .Z(state_7__N_911[5])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i14_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_192 (.A(n13141), .B(n87), .C(\PWMArray[0][9] ), 
         .D(n12221), .Z(\MATRIX_data[0] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(62[49:71])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_192.init = 16'h1000;
    LUT4 i2650_3_lut (.A(n5246), .B(n5245), .C(n5244), .Z(lastAddress_c[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(57[3] 106[10])
    defparam i2650_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PLL
//

module PLL (LOGIC_CLOCK_N_116, LOGIC_CLOCK, CLK_c, PIXEL_CLOCK, GND_net, 
            PIXEL_CLOCK_N_302) /* synthesis NGD_DRC_MASK=1 */ ;
    output LOGIC_CLOCK_N_116;
    output LOGIC_CLOCK;
    input CLK_c;
    output PIXEL_CLOCK;
    input GND_net;
    output PIXEL_CLOCK_N_302;
    
    wire LOGIC_CLOCK_N_116 /* synthesis is_clock=1, is_inv_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(73[9:17])
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire CLK_c /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(8[3:6])
    wire PIXEL_CLOCK /* synthesis SET_AS_NETWORK=PIXEL_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(43[8:19])
    wire PIXEL_CLOCK_N_302 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(82[9:22])
    
    INV i9642 (.A(LOGIC_CLOCK), .Z(LOGIC_CLOCK_N_116));
    EHXPLLJ PLLInst_0 (.CLKI(CLK_c), .CLKFB(LOGIC_CLOCK), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(LOGIC_CLOCK), .CLKOS(PIXEL_CLOCK)) /* synthesis FREQUENCY_PIN_CLKOS="35.416667", FREQUENCY_PIN_CLKOP="141.666667", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="8", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=13, LSE_LLINE=237, LSE_RLINE=237 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(237[10:13])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 17;
    defparam PLLInst_0.CLKOP_DIV = 4;
    defparam PLLInst_0.CLKOS_DIV = 16;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 3;
    defparam PLLInst_0.CLKOS_CPHASE = 15;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    INV i9643 (.A(PIXEL_CLOCK), .Z(PIXEL_CLOCK_N_302));
    
endmodule
//
// Verilog Description of module MatrixBusHandler
//

module MatrixBusHandler (\BUS_currGrantID[1] , \BUS_currGrantID[0] , \BUS_ADDR_INTERNAL[13] , 
            n13155, \BUS_ADDR_INTERNAL[14] , n13157, \BUS_ADDR_INTERNAL[11] , 
            n13156, \BUS_ADDR_INTERNAL[12] , n13142, n12248, n13158, 
            n12247, n1627, GND_net, \BUS_ADDR_INTERNAL[10] , n13143, 
            MATRIX_CURRROW, yOffset, n12342, LOGIC_CLOCK, n13160, 
            LOGIC_CLOCK_enable_71, BUS_data, \BUS_currGrantID_3__N_72[0] , 
            \VRAM_ADDR[0] , currReadRow, n12311, n12284, n12253, n12264, 
            n12259, n3116, n3117, n3118, n3119, n3112, n3113, 
            n3114, n3115, VRAM_WC, \BUS_ADDR_INTERNAL[0] , LOGIC_CLOCK_N_116, 
            n12219, n3132, n3133, n3134, n3135, n3217, n3218, 
            n3219, n3220, n3322, n3323, n3324, n3325, VRAM_DATA, 
            n12244, n10871, n3167, n3168, n3169, n3170, VCC_net, 
            n3027, \VRAM_ADDR[6] , \VRAM_ADDR[5] , \VRAM_ADDR[4] , MDM_done, 
            \VRAM_ADDR[3] , \VRAM_ADDR[2] , xOffset, \VRAM_ADDR[1] , 
            n3035, n3034, n3036, n3037, n3032, n3031, n3033, n3029, 
            n3028, n3030, LOGIC_CLOCK_enable_26, n5648, \BUS_ADDR_INTERNAL[18] , 
            \BUS_ADDR_INTERNAL[16] , \BUS_ADDR_INTERNAL[16]_adj_19 , \BUS_ADDR_INTERNAL[17] , 
            \lastReadRow[3] , \lastReadRow[4] , \BUS_ADDR_INTERNAL[15] , 
            \BUS_ADDR_INTERNAL[9] , \BUS_ADDR_INTERNAL[8] , \BUS_ADDR_INTERNAL[7] , 
            \BUS_ADDR_INTERNAL[6] , \BUS_ADDR_INTERNAL[5] , \BUS_ADDR_INTERNAL[4] , 
            \BUS_ADDR_INTERNAL[3] , \BUS_ADDR_INTERNAL[2] , \BUS_ADDR_INTERNAL[1] , 
            \BUS_ADDR_INTERNAL[14]_adj_20 , \BUS_ADDR_INTERNAL[15]_adj_21 , 
            \BUS_ADDR_INTERNAL[12]_adj_22 , \BUS_ADDR_INTERNAL[13]_adj_23 , 
            \otherData[7] , \BUS_DATA_INTERNAL[7] , \otherData[6] , \BUS_DATA_INTERNAL[6] , 
            \BUS_ADDR_INTERNAL[10]_adj_24 , \BUS_ADDR_INTERNAL[11]_adj_25 , 
            \otherData[5] , \BUS_DATA_INTERNAL[5] , \BUS_ADDR_INTERNAL[8]_adj_26 , 
            \BUS_ADDR_INTERNAL[9]_adj_27 , \otherData[4] , \BUS_DATA_INTERNAL[4] , 
            \BUS_ADDR_INTERNAL[6]_adj_28 , \BUS_ADDR_INTERNAL[7]_adj_29 , 
            \BUS_DATA_INTERNAL[3] , n3365, n3366, n3367, n3368, n3369, 
            n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3330, 
            n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
            n3339, n3340, n3341, n3349, n3350, n3351, n3352, n3353, 
            n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3314, 
            n3315, n3316, n3317, n3318, n3319, n3320, n3321, \BUS_DATA_INTERNAL[2] , 
            n3361, n3362, n3363, n3364, \BUS_DATA_INTERNAL[1] , \BUS_ADDR_INTERNAL[4]_adj_30 , 
            \BUS_ADDR_INTERNAL[5]_adj_31 , n3326, n3327, n3328, n3329, 
            n3342, n3343, n3344, n3345, \BUS_ADDR_INTERNAL[2]_adj_32 , 
            \BUS_ADDR_INTERNAL[3]_adj_33 , n3377, n3378, n3379, n3380, 
            n3260, n3261, n3262, n3263, n3278, n12277, n12344, 
            n12292, \BUS_DATA_INTERNAL[0] , n3264, n3265, n3266, n3267, 
            n3268, n3269, n3270, n3271, n3225, n3226, n3227, n3228, 
            n3243, n3229, n3230, n3231, n3232, n3233, n3234, n3235, 
            n3236, n3244, n3245, n3246, n3247, n3277, n3248, n3249, 
            n3250, n3251, n3252, n3253, n3254, n3255, n3209, n3210, 
            n3211, n3212, n12269, n3213, n3214, n3215, n3216, 
            n3256, n3257, n3258, n3259, n3221, n3222, n3223, n3224, 
            n3237, n3238, n3239, n3240, n3272, n3273, n3274, n3275, 
            n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
            n3163, n3164, n3165, n3166, n3120, n3121, n3122, n3123, 
            n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
            n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
            n3147, n3148, n3149, n3150, n3104, n3105, n3106, n3107, 
            n3108, n3109, n3110, n3111, n3151, n3152, n3153, n3154, 
            n12309, n13150, n13151, reset, n13144, n13154, LOGIC_CLOCK_enable_49, 
            n11094, n11095, n12263, n11096, n11097, n11150, n11151, 
            n11152, n11153, n11157, n11158, n11159, n11160, n11164, 
            n11165, n11166, n11167, n1921, n11171, n11172, n11174, 
            n11175, n11177, n11178, n11180, n11181, n11183, n11184, 
            n13146, n13147, n13153, n13145, n13152, n13148, n11101, 
            n11102, n13139, n12299, n11103, n11104, n12265, \MDM_data[13] , 
            \MDM_data[14] , n12261, n100, \BUS_DATA_INTERNAL[15] , n12218, 
            n4537, BUS_DONE, n11186, n11187, n4541, n63, n1184, 
            BUS_DONE_OUT_N_626, n4545, \MDM_data[8] , n11188, n11189, 
            \MDM_data[9] , n11193, n11194, \MDM_data[10] , n12329, 
            \MDM_data[11] , n13141, n12215, n11196, n11197, n12332, 
            n12352, n12222, n11199, n11200, \BUS_ADDR_INTERNAL[18]_derived_1 , 
            \MDM_data[12] , n11201, n11202, n11206, n11207, n11209, 
            n11210, n11212, n11213, n11215, n11216, n11217, n11218, 
            n12304, \lastAddress[18] , SRAM_WE_N_704, n46, n2025, 
            n13140, lastAddress_31__N_789, n12272, \BUS_addr[13] , lastAddress_31__N_845, 
            lastAddress_31__N_785, n12288, lastAddress_31__N_863, n12287, 
            lastAddress_31__N_787, lastAddress_31__N_783, n11222, n11223, 
            \BUS_addr[11] , lastAddress_31__N_779, lastAddress_31__N_851, 
            lastAddress_31__N_869, lastAddress_31__N_875, n12278, lastAddress_31__N_881, 
            lastAddress_31__N_777, \BUS_addr[14] , lastAddress_31__N_842, 
            lastAddress_31__N_776, n12291, lastAddress_31__N_857, lastAddress_31__N_872, 
            lastAddress_31__N_786, n11225, n11226, n11228, n11229, 
            n11231, n11232, n11234, n11235, n11237, n11238, n11108, 
            n11109, n11110, n11111, n11115, n11116, n12276, n11012, 
            n12274, n12273, n11117, n11118, n11122, n11123, n10350, 
            n10349, n11124, n11125, n11129, n11130, n11131, n11132, 
            n12280, n11324, n11325, n2266, n11326, n11327, n11136, 
            n11137, n10855, \lastAddress[1] , n63_adj_34, n2265, n11331, 
            n11332, n2264, n2263, n11333, n11334, n11138, n11139, 
            n11143, n11144, n11145, n11146, n12220, WRITE_DONE, 
            WRITE_DONE_adj_35, n7, BUS_DONE_OVERRIDE, BUS_DONE_INTERNAL, 
            \GR_WR_ADDR[6] , \GR_WR_ADDR[2] , \GR_WR_ADDR[0] , \GR_WR_DOUT[7] , 
            \GR_WR_DOUT[6] , \GR_WR_DOUT[5] , \GR_WR_DOUT[4] );
    input \BUS_currGrantID[1] ;
    input \BUS_currGrantID[0] ;
    output \BUS_ADDR_INTERNAL[13] ;
    input n13155;
    output \BUS_ADDR_INTERNAL[14] ;
    input n13157;
    output \BUS_ADDR_INTERNAL[11] ;
    input n13156;
    output \BUS_ADDR_INTERNAL[12] ;
    input n13142;
    input n12248;
    output n13158;
    input n12247;
    output n1627;
    input GND_net;
    output \BUS_ADDR_INTERNAL[10] ;
    input n13143;
    input [4:0]MATRIX_CURRROW;
    output [7:0]yOffset;
    input n12342;
    input LOGIC_CLOCK;
    input n13160;
    input LOGIC_CLOCK_enable_71;
    output [15:0]BUS_data;
    output \BUS_currGrantID_3__N_72[0] ;
    output \VRAM_ADDR[0] ;
    input [4:0]currReadRow;
    input n12311;
    input n12284;
    input n12253;
    input n12264;
    input n12259;
    output n3116;
    output n3117;
    output n3118;
    output n3119;
    output n3112;
    output n3113;
    output n3114;
    output n3115;
    output VRAM_WC;
    output \BUS_ADDR_INTERNAL[0] ;
    input LOGIC_CLOCK_N_116;
    output n12219;
    output n3132;
    output n3133;
    output n3134;
    output n3135;
    output n3217;
    output n3218;
    output n3219;
    output n3220;
    output n3322;
    output n3323;
    output n3324;
    output n3325;
    output [9:0]VRAM_DATA;
    input n12244;
    input n10871;
    output n3167;
    output n3168;
    output n3169;
    output n3170;
    input VCC_net;
    output [9:0]n3027;
    output \VRAM_ADDR[6] ;
    output \VRAM_ADDR[5] ;
    output \VRAM_ADDR[4] ;
    output MDM_done;
    output \VRAM_ADDR[3] ;
    output \VRAM_ADDR[2] ;
    output [7:0]xOffset;
    output \VRAM_ADDR[1] ;
    output [9:0]n3035;
    output [9:0]n3034;
    output [9:0]n3036;
    output [9:0]n3037;
    output [9:0]n3032;
    output [9:0]n3031;
    output [9:0]n3033;
    output [9:0]n3029;
    output [9:0]n3028;
    output [9:0]n3030;
    input LOGIC_CLOCK_enable_26;
    input n5648;
    input \BUS_ADDR_INTERNAL[18] ;
    input \BUS_ADDR_INTERNAL[16] ;
    output \BUS_ADDR_INTERNAL[16]_adj_19 ;
    input \BUS_ADDR_INTERNAL[17] ;
    output \lastReadRow[3] ;
    output \lastReadRow[4] ;
    output \BUS_ADDR_INTERNAL[15] ;
    output \BUS_ADDR_INTERNAL[9] ;
    output \BUS_ADDR_INTERNAL[8] ;
    output \BUS_ADDR_INTERNAL[7] ;
    output \BUS_ADDR_INTERNAL[6] ;
    output \BUS_ADDR_INTERNAL[5] ;
    output \BUS_ADDR_INTERNAL[4] ;
    output \BUS_ADDR_INTERNAL[3] ;
    output \BUS_ADDR_INTERNAL[2] ;
    output \BUS_ADDR_INTERNAL[1] ;
    input \BUS_ADDR_INTERNAL[14]_adj_20 ;
    input \BUS_ADDR_INTERNAL[15]_adj_21 ;
    input \BUS_ADDR_INTERNAL[12]_adj_22 ;
    input \BUS_ADDR_INTERNAL[13]_adj_23 ;
    input \otherData[7] ;
    output \BUS_DATA_INTERNAL[7] ;
    input \otherData[6] ;
    output \BUS_DATA_INTERNAL[6] ;
    input \BUS_ADDR_INTERNAL[10]_adj_24 ;
    input \BUS_ADDR_INTERNAL[11]_adj_25 ;
    input \otherData[5] ;
    output \BUS_DATA_INTERNAL[5] ;
    input \BUS_ADDR_INTERNAL[8]_adj_26 ;
    input \BUS_ADDR_INTERNAL[9]_adj_27 ;
    input \otherData[4] ;
    output \BUS_DATA_INTERNAL[4] ;
    input \BUS_ADDR_INTERNAL[6]_adj_28 ;
    input \BUS_ADDR_INTERNAL[7]_adj_29 ;
    output \BUS_DATA_INTERNAL[3] ;
    output n3365;
    output n3366;
    output n3367;
    output n3368;
    output n3369;
    output n3370;
    output n3371;
    output n3372;
    output n3373;
    output n3374;
    output n3375;
    output n3376;
    output n3330;
    output n3331;
    output n3332;
    output n3333;
    output n3334;
    output n3335;
    output n3336;
    output n3337;
    output n3338;
    output n3339;
    output n3340;
    output n3341;
    output n3349;
    output n3350;
    output n3351;
    output n3352;
    output n3353;
    output n3354;
    output n3355;
    output n3356;
    output n3357;
    output n3358;
    output n3359;
    output n3360;
    output n3314;
    output n3315;
    output n3316;
    output n3317;
    output n3318;
    output n3319;
    output n3320;
    output n3321;
    output \BUS_DATA_INTERNAL[2] ;
    output n3361;
    output n3362;
    output n3363;
    output n3364;
    output \BUS_DATA_INTERNAL[1] ;
    input \BUS_ADDR_INTERNAL[4]_adj_30 ;
    input \BUS_ADDR_INTERNAL[5]_adj_31 ;
    output n3326;
    output n3327;
    output n3328;
    output n3329;
    output n3342;
    output n3343;
    output n3344;
    output n3345;
    input \BUS_ADDR_INTERNAL[2]_adj_32 ;
    input \BUS_ADDR_INTERNAL[3]_adj_33 ;
    output n3377;
    output n3378;
    output n3379;
    output n3380;
    output n3260;
    output n3261;
    output n3262;
    output n3263;
    input n3278;
    input n12277;
    input n12344;
    input n12292;
    output \BUS_DATA_INTERNAL[0] ;
    output n3264;
    output n3265;
    output n3266;
    output n3267;
    output n3268;
    output n3269;
    output n3270;
    output n3271;
    output n3225;
    output n3226;
    output n3227;
    output n3228;
    input n3243;
    output n3229;
    output n3230;
    output n3231;
    output n3232;
    output n3233;
    output n3234;
    output n3235;
    output n3236;
    output n3244;
    output n3245;
    output n3246;
    output n3247;
    input n3277;
    output n3248;
    output n3249;
    output n3250;
    output n3251;
    output n3252;
    output n3253;
    output n3254;
    output n3255;
    output n3209;
    output n3210;
    output n3211;
    output n3212;
    input n12269;
    output n3213;
    output n3214;
    output n3215;
    output n3216;
    output n3256;
    output n3257;
    output n3258;
    output n3259;
    output n3221;
    output n3222;
    output n3223;
    output n3224;
    output n3237;
    output n3238;
    output n3239;
    output n3240;
    output n3272;
    output n3273;
    output n3274;
    output n3275;
    output n3155;
    output n3156;
    output n3157;
    output n3158;
    output n3159;
    output n3160;
    output n3161;
    output n3162;
    output n3163;
    output n3164;
    output n3165;
    output n3166;
    output n3120;
    output n3121;
    output n3122;
    output n3123;
    output n3124;
    output n3125;
    output n3126;
    output n3127;
    output n3128;
    output n3129;
    output n3130;
    output n3131;
    output n3139;
    output n3140;
    output n3141;
    output n3142;
    output n3143;
    output n3144;
    output n3145;
    output n3146;
    output n3147;
    output n3148;
    output n3149;
    output n3150;
    output n3104;
    output n3105;
    output n3106;
    output n3107;
    output n3108;
    output n3109;
    output n3110;
    output n3111;
    output n3151;
    output n3152;
    output n3153;
    output n3154;
    input n12309;
    input n13150;
    input n13151;
    output reset;
    input n13144;
    input n13154;
    input LOGIC_CLOCK_enable_49;
    input n11094;
    input n11095;
    input n12263;
    input n11096;
    input n11097;
    input n11150;
    input n11151;
    input n11152;
    input n11153;
    input n11157;
    input n11158;
    input n11159;
    input n11160;
    input n11164;
    input n11165;
    input n11166;
    input n11167;
    output n1921;
    input n11171;
    input n11172;
    input n11174;
    input n11175;
    input n11177;
    input n11178;
    input n11180;
    input n11181;
    input n11183;
    input n11184;
    input n13146;
    input n13147;
    input n13153;
    input n13145;
    input n13152;
    input n13148;
    input n11101;
    input n11102;
    input n13139;
    input n12299;
    input n11103;
    input n11104;
    input n12265;
    output \MDM_data[13] ;
    output \MDM_data[14] ;
    input n12261;
    input n100;
    input \BUS_DATA_INTERNAL[15] ;
    output n12218;
    input n4537;
    output BUS_DONE;
    input n11186;
    input n11187;
    input n4541;
    input n63;
    input n1184;
    input BUS_DONE_OUT_N_626;
    input n4545;
    output \MDM_data[8] ;
    input n11188;
    input n11189;
    output \MDM_data[9] ;
    input n11193;
    input n11194;
    output \MDM_data[10] ;
    output n12329;
    output \MDM_data[11] ;
    input n13141;
    output n12215;
    input n11196;
    input n11197;
    input n12332;
    input n12352;
    input n12222;
    input n11199;
    input n11200;
    input \BUS_ADDR_INTERNAL[18]_derived_1 ;
    output \MDM_data[12] ;
    input n11201;
    input n11202;
    input n11206;
    input n11207;
    input n11209;
    input n11210;
    input n11212;
    input n11213;
    input n11215;
    input n11216;
    input n11217;
    input n11218;
    input n12304;
    input \lastAddress[18] ;
    input SRAM_WE_N_704;
    output n46;
    output n2025;
    input n13140;
    output lastAddress_31__N_789;
    input n12272;
    input \BUS_addr[13] ;
    output lastAddress_31__N_845;
    output lastAddress_31__N_785;
    input n12288;
    output lastAddress_31__N_863;
    input n12287;
    output lastAddress_31__N_787;
    output lastAddress_31__N_783;
    input n11222;
    input n11223;
    input \BUS_addr[11] ;
    output lastAddress_31__N_779;
    output lastAddress_31__N_851;
    output lastAddress_31__N_869;
    output lastAddress_31__N_875;
    input n12278;
    output lastAddress_31__N_881;
    output lastAddress_31__N_777;
    input \BUS_addr[14] ;
    output lastAddress_31__N_842;
    output lastAddress_31__N_776;
    input n12291;
    output lastAddress_31__N_857;
    output lastAddress_31__N_872;
    output lastAddress_31__N_786;
    input n11225;
    input n11226;
    input n11228;
    input n11229;
    input n11231;
    input n11232;
    input n11234;
    input n11235;
    input n11237;
    input n11238;
    input n11108;
    input n11109;
    input n11110;
    input n11111;
    input n11115;
    input n11116;
    input n12276;
    input n11012;
    input n12274;
    input n12273;
    input n11117;
    input n11118;
    input n11122;
    input n11123;
    input n10350;
    input n10349;
    input n11124;
    input n11125;
    input n11129;
    input n11130;
    input n11131;
    input n11132;
    input n12280;
    input n11324;
    input n11325;
    input n2266;
    input n11326;
    input n11327;
    input n11136;
    input n11137;
    input n10855;
    input \lastAddress[1] ;
    output n63_adj_34;
    input n2265;
    input n11331;
    input n11332;
    input n2264;
    input n2263;
    input n11333;
    input n11334;
    input n11138;
    input n11139;
    input n11143;
    input n11144;
    input n11145;
    input n11146;
    input n12220;
    input WRITE_DONE;
    input WRITE_DONE_adj_35;
    input n7;
    input BUS_DONE_OVERRIDE;
    input BUS_DONE_INTERNAL;
    input \GR_WR_ADDR[6] ;
    input \GR_WR_ADDR[2] ;
    input \GR_WR_ADDR[0] ;
    output \GR_WR_DOUT[7] ;
    output \GR_WR_DOUT[6] ;
    output \GR_WR_DOUT[5] ;
    output \GR_WR_DOUT[4] ;
    
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire MATRIX_CURRROW_0_derived_5 /* synthesis is_clock=1, SET_AS_NETWORK=MATRIX_CURRROW[0]_derived_5 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(91[8:22])
    wire offsetLatchClockOrd /* synthesis is_clock=1, SET_AS_NETWORK=\MDM/offsetLatchClockOrd */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(59[9:28])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(90[8:15])
    wire LOGIC_CLOCK_N_116 /* synthesis is_clock=1, is_inv_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(73[9:17])
    wire GR_WR_CLK /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(138[9:18])
    
    wire n10200, n10201, n10199, n12, n9981;
    wire [7:0]y;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(68[9:10])
    
    wire n9982, frameEndClock, LOGIC_CLOCK_enable_1;
    wire [7:0]xOffset_pre;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(60[9:20])
    
    wire LOGIC_CLOCK_enable_6, n10852;
    wire [7:0]yOffset_pre;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(61[9:20])
    
    wire n12232;
    wire [1:0]currRowOffset_lat;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(77[9:26])
    
    wire n3291;
    wire [7:0]state;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    
    wire n10478, LOGIC_CLOCK_enable_175;
    wire [8:0]n280;
    wire [4:0]lastReadRow;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(55[9:20])
    
    wire n9983, n3137;
    wire [1:0]currRowOffset;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(74[9:22])
    
    wire VRAM_WC_N_598;
    wire [3:0]currColor_lat;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(78[9:22])
    wire [3:0]currColor;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(72[9:18])
    
    wire LOGIC_CLOCK_N_116_enable_20;
    wire [31:0]currAddress;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(73[9:20])
    wire [3:0]BUS_transferState;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(109[9:26])
    
    wire LOGIC_CLOCK_enable_10, n3138, n3242, n3347;
    wire [9:0]GR_RE_DOUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(135[9:19])
    
    wire n3296, n10898, LOGIC_CLOCK_enable_78, n3173;
    wire [3:0]latchMode;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(121[9:18])
    
    wire LOGIC_CLOCK_enable_81, LOGIC_CLOCK_enable_16, n3306, n3301;
    wire [17:0]currAddress_17__N_488;
    
    wire n10166, n1956, GR_WR_CLK_N_689, n10165, n10164;
    wire [31:0]BUS_ADDR_INTERNAL;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(81[9:26])
    wire [7:0]xPre;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(69[9:13])
    
    wire LOGIC_CLOCK_enable_167;
    wire [7:0]n37;
    
    wire n14, n54, n24, n10163, n10162;
    wire [15:0]Sprite_readData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(95[9:24])
    
    wire n11093, n10161;
    wire [1:0]n1;
    
    wire n10436, n10160, n10870, n10159;
    wire [15:0]otherData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(97[9:18])
    wire [7:0]n2372;
    
    wire n10540, n3383, n3348, n3382, n9979;
    wire [7:0]x;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(67[9:10])
    
    wire n10158, n10157, n9978, n11147, n11148, n11149, n11154, 
        n11155, n11156, n11098, n11099, n11100, n12049, n11161, 
        n11162, n11163, n11168, n11169, n11170, n11105, n11106, 
        n11107, n3172, n11190, n11191, n11192, n10136, n2129, 
        n11203, n11204, n11205;
    wire [7:0]currValue;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(75[9:18])
    
    wire LOGIC_CLOCK_enable_178;
    wire [3:0]n27;
    
    wire n10135, n11219, n11220, n11221, n10134, n10133, state_7__N_322, 
        reset_N_670, n11112, n11113, n11114, n10132, n10131, n10130, 
        latchForce, n11119, n11120, n11121, n11126, n11127, n11128, 
        n11133, n11134, n11135, n11328, n11329, n11330, n11335, 
        n11336, n11337, n11140, n11141, n11142, n10084, n9977;
    wire [15:0]Sprite_readData_15__N_417;
    
    wire n10083, n10082, n10081, n10080, n10079, n9995;
    wire [9:0]currAddress_17__N_506;
    
    wire n10078, n9994, n10077, n10076, n10075, n9993, n9992, 
        n10309, n13, n12331, BUS_DONE_OUT_N_627, n12230, n10846, 
        BUS_VALID_N_480, n3790;
    wire [9:0]GR_WR_DOUT;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(133[9:19])
    
    wire n10042, n10041, n4, n10348, n12092, n10040, n4_adj_1294;
    wire [7:0]n162;
    
    wire n9984, n10039, n12226, n8, n12228, n12_adj_1295, n12224, 
        n18, n11052, n12157, n12050, n12048, n10033, n10032;
    wire [7:0]GR_WR_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(136[9:19])
    
    wire n10031, n10030, n12343, n10029, n13_adj_1297, n11, n15_adj_1298, 
        n8148, n10028, n10027, n12338, n11068, n8_adj_1299, n6, 
        n12327, n19, n160, n10026, n10025, n10024, n12297, n11_adj_1301, 
        n10023, n10893, n9, n10022, n21, n10021, n10204, n10203, 
        n11060, n10202, n10888, n10;
    
    CCU2D add_7182_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n13155), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n13157), 
          .CIN(n10200), .COUT(n10201));
    defparam add_7182_5.INIT0 = 16'h00ae;
    defparam add_7182_5.INIT1 = 16'h00ae;
    defparam add_7182_5.INJECT1_0 = "NO";
    defparam add_7182_5.INJECT1_1 = "NO";
    CCU2D add_7182_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n13156), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n13142), 
          .CIN(n10199), .COUT(n10200));
    defparam add_7182_3.INIT0 = 16'h00ae;
    defparam add_7182_3.INIT1 = 16'h00ae;
    defparam add_7182_3.INJECT1_0 = "NO";
    defparam add_7182_3.INJECT1_1 = "NO";
    LUT4 i6_4_lut (.A(n12248), .B(n12), .C(n13158), .D(n12247), .Z(n1627)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i6_4_lut.init = 16'h0080;
    CCU2D add_7182_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), 
          .D1(n13143), .COUT(n10199));
    defparam add_7182_1.INIT0 = 16'hF000;
    defparam add_7182_1.INIT1 = 16'h00ae;
    defparam add_7182_1.INJECT1_0 = "NO";
    defparam add_7182_1.INJECT1_1 = "NO";
    CCU2D yPre_7__I_0_3 (.A0(MATRIX_CURRROW[1]), .B0(MATRIX_CURRROW[0]), 
          .C0(yOffset[1]), .D0(GND_net), .A1(MATRIX_CURRROW[2]), .B1(n12342), 
          .C1(yOffset[2]), .D1(GND_net), .CIN(n9981), .COUT(n9982), 
          .S0(y[1]), .S1(y[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(165[24:38])
    defparam yPre_7__I_0_3.INIT0 = 16'h9696;
    defparam yPre_7__I_0_3.INIT1 = 16'h9696;
    defparam yPre_7__I_0_3.INJECT1_0 = "NO";
    defparam yPre_7__I_0_3.INJECT1_1 = "NO";
    FD1P3DX frameEndClock_343 (.D(n13160), .SP(LOGIC_CLOCK_enable_1), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(frameEndClock)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam frameEndClock_343.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i0.GSR = "DISABLED";
    FD1P3AX BUS_REQ_345 (.D(n10852), .SP(LOGIC_CLOCK_enable_6), .CK(LOGIC_CLOCK), 
            .Q(\BUS_currGrantID_3__N_72[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam BUS_REQ_345.GSR = "DISABLED";
    FD1S3AX yOffset_i0 (.D(yOffset_pre[0]), .CK(offsetLatchClockOrd), .Q(yOffset[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(n12232), .B(currRowOffset_lat[0]), .C(currRowOffset_lat[1]), 
         .Z(n3291)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0202;
    FD1S3DX state__i0 (.D(n10478), .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), 
            .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam state__i0.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i1 (.D(n280[0]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i1.GSR = "DISABLED";
    FD1S1A currReadRow_4__I_0_424_i1 (.D(currReadRow[0]), .CK(MATRIX_CURRROW_0_derived_5), 
           .Q(lastReadRow[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[2] 275[14])
    defparam currReadRow_4__I_0_424_i1.GSR = "DISABLED";
    CCU2D yPre_7__I_0_5 (.A0(MATRIX_CURRROW[3]), .B0(n12311), .C0(yOffset[3]), 
          .D0(GND_net), .A1(MATRIX_CURRROW[4]), .B1(n12284), .C1(yOffset[4]), 
          .D1(GND_net), .CIN(n9982), .COUT(n9983), .S0(y[3]), .S1(y[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(165[24:38])
    defparam yPre_7__I_0_5.INIT0 = 16'h9696;
    defparam yPre_7__I_0_5.INIT1 = 16'h9696;
    defparam yPre_7__I_0_5.INJECT1_0 = "NO";
    defparam yPre_7__I_0_5.INJECT1_1 = "NO";
    SPR16X4C Sprite_positions3 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), 
            .AD2(n12259), .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3137), 
            .DO0(n3116), .DO1(n3117), .DO2(n3118), .DO3(n3119));
    defparam Sprite_positions3.initval = "0x0000000000000000";
    FD1P3AX currRowOffset_lat_i0_i0 (.D(currRowOffset[0]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currRowOffset_lat[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currRowOffset_lat_i0_i0.GSR = "DISABLED";
    SPR16X4C Sprite_positions4 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3137), .DO0(n3112), 
            .DO1(n3113), .DO2(n3114), .DO3(n3115));
    defparam Sprite_positions4.initval = "0x0000000000000000";
    FD1S3DX VRAM_WC_339 (.D(VRAM_WC_N_598), .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), 
            .Q(VRAM_WC)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_WC_339.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i0 (.D(currColor[0]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currColor_lat_i0_i0.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i1 (.D(currAddress[0]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i1.GSR = "DISABLED";
    FD1P3DX BUS_transferState__i1 (.D(n13160), .SP(LOGIC_CLOCK_enable_10), 
            .CK(LOGIC_CLOCK), .CD(n12219), .Q(BUS_transferState[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam BUS_transferState__i1.GSR = "DISABLED";
    SPR16X4C Sprite_positions1 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), 
            .AD2(n12259), .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3138), 
            .DO0(n3132), .DO1(n3133), .DO2(n3134), .DO3(n3135));
    defparam Sprite_positions1.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes4 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3242), .DO0(n3217), 
            .DO1(n3218), .DO2(n3219), .DO3(n3220));
    defparam Sprite_sizes4.initval = "0x0000000000000000";
    SPR16X4C Sprite_options4 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3347), .DO0(n3322), 
            .DO1(n3323), .DO2(n3324), .DO3(n3325));
    defparam Sprite_options4.initval = "0x0000000000000000";
    DPR16X4C n30401 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(VRAM_DATA[2]), .DO1(VRAM_DATA[3]), .DO2(VRAM_DATA[4]), 
            .DO3(VRAM_DATA[5]));
    defparam n30401.initval = "0x0000000000000000";
    LUT4 i5_4_lut (.A(n12264), .B(n12244), .C(n10871), .D(n10898), .Z(n12)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i5_4_lut.init = 16'h1000;
    FD1P3AX yOffset_pre_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i0.GSR = "DISABLED";
    SPR16X4C Sprite_positions2 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), 
            .AD2(n12259), .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3173), 
            .DO0(n3167), .DO1(n3168), .DO2(n3169), .DO3(n3170));
    defparam Sprite_positions2.initval = "0x0000000000000000";
    DPR16X4C n3039_d02 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3027[0]), .DO1(n3027[1]));
    defparam n3039_d02.initval = "0x0000000000000000";
    FD1P3AX latchMode_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_81), 
            .CK(LOGIC_CLOCK), .Q(latchMode[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam latchMode_i0_i0.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i7 (.D(n280[6]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i7.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i6 (.D(n280[5]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i6.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i5 (.D(n280[4]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i5.GSR = "DISABLED";
    FD1P3DX transferDone_363 (.D(n13160), .SP(LOGIC_CLOCK_enable_16), .CK(LOGIC_CLOCK), 
            .CD(n12219), .Q(MDM_done)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam transferDone_363.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i4 (.D(n280[3]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i4.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i3 (.D(n280[2]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i3.GSR = "DISABLED";
    FD1S3AX xOffset_i0 (.D(xOffset_pre[0]), .CK(offsetLatchClockOrd), .Q(xOffset[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i0.GSR = "DISABLED";
    FD1P3AX VRAM_ADDR__i2 (.D(n280[1]), .SP(LOGIC_CLOCK_enable_175), .CK(LOGIC_CLOCK), 
            .Q(\VRAM_ADDR[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam VRAM_ADDR__i2.GSR = "DISABLED";
    DPR16X4C n30461 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3035[2]), .DO1(n3035[3]), .DO2(n3035[4]), .DO3(n3035[5]));
    defparam n30461.initval = "0x0000000000000000";
    DPR16X4C n3044_d51 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3034[2]), .DO1(n3034[3]), .DO2(n3034[4]), .DO3(n3034[5]));
    defparam n3044_d51.initval = "0x0000000000000000";
    DPR16X4C n3045_d61 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3036[2]), .DO1(n3036[3]), .DO2(n3036[4]), .DO3(n3036[5]));
    defparam n3045_d61.initval = "0x0000000000000000";
    DPR16X4C n3039_d01 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3027[2]), .DO1(n3027[3]), .DO2(n3027[4]), .DO3(n3027[5]));
    defparam n3039_d01.initval = "0x0000000000000000";
    DPR16X4C n3046_d71 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3037[2]), .DO1(n3037[3]), .DO2(n3037[4]), .DO3(n3037[5]));
    defparam n3046_d71.initval = "0x0000000000000000";
    DPR16X4C n30441 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3032[2]), .DO1(n3032[3]), .DO2(n3032[4]), .DO3(n3032[5]));
    defparam n30441.initval = "0x0000000000000000";
    DPR16X4C n3042_d31 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3031[2]), .DO1(n3031[3]), .DO2(n3031[4]), .DO3(n3031[5]));
    defparam n3042_d31.initval = "0x0000000000000000";
    DPR16X4C n3043_d41 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3033[2]), .DO1(n3033[3]), .DO2(n3033[4]), .DO3(n3033[5]));
    defparam n3043_d41.initval = "0x0000000000000000";
    DPR16X4C n30421 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3029[2]), .DO1(n3029[3]), .DO2(n3029[4]), .DO3(n3029[5]));
    defparam n30421.initval = "0x0000000000000000";
    DPR16X4C n3040_d11 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3028[2]), .DO1(n3028[3]), .DO2(n3028[4]), .DO3(n3028[5]));
    defparam n3040_d11.initval = "0x0000000000000000";
    DPR16X4C n3041_d21 (.DI0(GR_RE_DOUT[2]), .DI1(GR_RE_DOUT[3]), .DI2(GR_RE_DOUT[4]), 
            .DI3(GR_RE_DOUT[5]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3030[2]), .DO1(n3030[3]), .DO2(n3030[4]), .DO3(n3030[5]));
    defparam n3041_d21.initval = "0x0000000000000000";
    DPR16X4C n3041_d22 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3030[0]), .DO1(n3030[1]));
    defparam n3041_d22.initval = "0x0000000000000000";
    DPR16X4C n3040_d12 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3028[0]), .DO1(n3028[1]));
    defparam n3040_d12.initval = "0x0000000000000000";
    DPR16X4C n3042_d32 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3031[0]), .DO1(n3031[1]));
    defparam n3042_d32.initval = "0x0000000000000000";
    DPR16X4C n3043_d42 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3033[0]), .DO1(n3033[1]));
    defparam n3043_d42.initval = "0x0000000000000000";
    LUT4 i1_2_lut_3_lut_adj_148 (.A(n12232), .B(currRowOffset_lat[0]), .C(currRowOffset_lat[1]), 
         .Z(n3296)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_148.init = 16'h0808;
    CCU2D yPre_7__I_0_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(MATRIX_CURRROW[0]), .B1(yOffset[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n9981), .S1(currAddress_17__N_488[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(165[24:38])
    defparam yPre_7__I_0_1.INIT0 = 16'hF000;
    defparam yPre_7__I_0_1.INIT1 = 16'ha999;
    defparam yPre_7__I_0_1.INJECT1_0 = "NO";
    defparam yPre_7__I_0_1.INJECT1_1 = "NO";
    CCU2D add_7184_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10166), .S1(n1956));
    defparam add_7184_21.INIT0 = 16'h1eee;
    defparam add_7184_21.INIT1 = 16'h0000;
    defparam add_7184_21.INJECT1_0 = "NO";
    defparam add_7184_21.INJECT1_1 = "NO";
    FD1P3DX GR_WR_CLK_364 (.D(GR_WR_CLK_N_689), .SP(LOGIC_CLOCK_enable_26), 
            .CK(LOGIC_CLOCK), .CD(n12219), .Q(GR_WR_CLK)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam GR_WR_CLK_364.GSR = "DISABLED";
    DPR16X4C n3045_d62 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3036[0]), .DO1(n3036[1]));
    defparam n3045_d62.initval = "0x0000000000000000";
    CCU2D add_7184_19 (.A0(n5648), .B0(\BUS_currGrantID[1] ), .C0(\BUS_currGrantID[0] ), 
          .D0(\BUS_ADDR_INTERNAL[18] ), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n10165), .COUT(n10166));
    defparam add_7184_19.INIT0 = 16'h0703;
    defparam add_7184_19.INIT1 = 16'h1eee;
    defparam add_7184_19.INJECT1_0 = "NO";
    defparam add_7184_19.INJECT1_1 = "NO";
    CCU2D add_7184_17 (.A0(\BUS_ADDR_INTERNAL[16] ), .B0(\BUS_ADDR_INTERNAL[16]_adj_19 ), 
          .C0(\BUS_currGrantID[0] ), .D0(\BUS_currGrantID[1] ), .A1(BUS_ADDR_INTERNAL[17]), 
          .B1(\BUS_ADDR_INTERNAL[17] ), .C1(\BUS_currGrantID[1] ), .D1(\BUS_currGrantID[0] ), 
          .CIN(n10164), .COUT(n10165));
    defparam add_7184_17.INIT0 = 16'h0acf;
    defparam add_7184_17.INIT1 = 16'hf530;
    defparam add_7184_17.INJECT1_0 = "NO";
    defparam add_7184_17.INJECT1_1 = "NO";
    DPR16X4C n3046_d72 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3037[0]), .DO1(n3037[1]));
    defparam n3046_d72.initval = "0x0000000000000000";
    FD1S1A currReadRow_4__I_0_424_i2 (.D(currReadRow[1]), .CK(MATRIX_CURRROW_0_derived_5), 
           .Q(lastReadRow[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[2] 275[14])
    defparam currReadRow_4__I_0_424_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_149 (.A(n12232), .B(currRowOffset_lat[0]), .C(currRowOffset_lat[1]), 
         .Z(n3306)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_149.init = 16'h8080;
    FD1S1A currReadRow_4__I_0_424_i3 (.D(currReadRow[2]), .CK(MATRIX_CURRROW_0_derived_5), 
           .Q(lastReadRow[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[2] 275[14])
    defparam currReadRow_4__I_0_424_i3.GSR = "DISABLED";
    FD1S1A currReadRow_4__I_0_424_i4 (.D(currReadRow[3]), .CK(MATRIX_CURRROW_0_derived_5), 
           .Q(\lastReadRow[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[2] 275[14])
    defparam currReadRow_4__I_0_424_i4.GSR = "DISABLED";
    FD1S1A currReadRow_4__I_0_424_i5 (.D(currReadRow[4]), .CK(MATRIX_CURRROW_0_derived_5), 
           .Q(\lastReadRow[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(182[2] 275[14])
    defparam currReadRow_4__I_0_424_i5.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i18 (.D(currAddress[17]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(BUS_ADDR_INTERNAL[17])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i18.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i17 (.D(currAddress[16]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[16]_adj_19 )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i17.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i16 (.D(currAddress[15]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[15] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i16.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i15 (.D(currAddress[14]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[14] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i15.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i14 (.D(currAddress[13]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[13] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i14.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i13 (.D(currAddress[12]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i13.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i12 (.D(currAddress[11]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i12.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i11 (.D(currAddress[10]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i11.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i10 (.D(currAddress[9]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i10.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i9 (.D(currAddress[8]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i9.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i8 (.D(currAddress[7]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i8.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i7 (.D(currAddress[6]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i7.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i6 (.D(currAddress[5]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i6.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i5 (.D(currAddress[4]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i5.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i4 (.D(currAddress[3]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i4.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i3 (.D(currAddress[2]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i3.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i2 (.D(currAddress[1]), .SP(LOGIC_CLOCK_N_116_enable_20), 
            .CK(LOGIC_CLOCK_N_116), .Q(\BUS_ADDR_INTERNAL[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(270[3] 274[10])
    defparam BUS_ADDR_INTERNAL__i2.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i3 (.D(currColor[3]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currColor_lat_i0_i3.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i2 (.D(currColor[2]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currColor_lat_i0_i2.GSR = "DISABLED";
    FD1P3AX currColor_lat_i0_i1 (.D(currColor[1]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currColor_lat[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currColor_lat_i0_i1.GSR = "DISABLED";
    FD1P3AX currRowOffset_lat_i0_i1 (.D(currRowOffset[1]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currRowOffset_lat[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currRowOffset_lat_i0_i1.GSR = "DISABLED";
    FD1P3DX xPre_681__i0 (.D(n37[0]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[0])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i0.GSR = "DISABLED";
    PFUMX i41 (.BLUT(n14), .ALUT(n54), .C0(state[0]), .Z(n24));
    CCU2D add_7184_15 (.A0(\BUS_ADDR_INTERNAL[14]_adj_20 ), .B0(\BUS_ADDR_INTERNAL[14] ), 
          .C0(\BUS_currGrantID[0] ), .D0(\BUS_currGrantID[1] ), .A1(\BUS_ADDR_INTERNAL[15]_adj_21 ), 
          .B1(\BUS_ADDR_INTERNAL[15] ), .C1(\BUS_currGrantID[0] ), .D1(\BUS_currGrantID[1] ), 
          .CIN(n10163), .COUT(n10164));
    defparam add_7184_15.INIT0 = 16'hf530;
    defparam add_7184_15.INIT1 = 16'hf530;
    defparam add_7184_15.INJECT1_0 = "NO";
    defparam add_7184_15.INJECT1_1 = "NO";
    CCU2D add_7184_13 (.A0(\BUS_ADDR_INTERNAL[12]_adj_22 ), .B0(\BUS_ADDR_INTERNAL[12] ), 
          .C0(\BUS_currGrantID[0] ), .D0(\BUS_currGrantID[1] ), .A1(\BUS_ADDR_INTERNAL[13]_adj_23 ), 
          .B1(\BUS_ADDR_INTERNAL[13] ), .C1(\BUS_currGrantID[0] ), .D1(\BUS_currGrantID[1] ), 
          .CIN(n10162), .COUT(n10163));
    defparam add_7184_13.INIT0 = 16'hf530;
    defparam add_7184_13.INIT1 = 16'hf530;
    defparam add_7184_13.INJECT1_0 = "NO";
    defparam add_7184_13.INJECT1_1 = "NO";
    PFUMX mux_472_i8 (.BLUT(Sprite_readData[7]), .ALUT(\otherData[7] ), 
          .C0(n11093), .Z(\BUS_DATA_INTERNAL[7] ));
    PFUMX mux_472_i7 (.BLUT(Sprite_readData[6]), .ALUT(\otherData[6] ), 
          .C0(n11093), .Z(\BUS_DATA_INTERNAL[6] ));
    CCU2D add_7184_11 (.A0(\BUS_ADDR_INTERNAL[10]_adj_24 ), .B0(\BUS_ADDR_INTERNAL[10] ), 
          .C0(\BUS_currGrantID[0] ), .D0(\BUS_currGrantID[1] ), .A1(\BUS_ADDR_INTERNAL[11]_adj_25 ), 
          .B1(\BUS_ADDR_INTERNAL[11] ), .C1(\BUS_currGrantID[0] ), .D1(\BUS_currGrantID[1] ), 
          .CIN(n10161), .COUT(n10162));
    defparam add_7184_11.INIT0 = 16'hf530;
    defparam add_7184_11.INIT1 = 16'hf530;
    defparam add_7184_11.INJECT1_0 = "NO";
    defparam add_7184_11.INJECT1_1 = "NO";
    FD1P3DX currRowOffset_682__i0 (.D(n1[0]), .SP(LOGIC_CLOCK_enable_167), 
            .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), .Q(currRowOffset[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currRowOffset_682__i0.GSR = "DISABLED";
    FD1S3DX state__i4 (.D(n10436), .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), 
            .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam state__i4.GSR = "DISABLED";
    PFUMX mux_472_i6 (.BLUT(Sprite_readData[5]), .ALUT(\otherData[5] ), 
          .C0(n11093), .Z(\BUS_DATA_INTERNAL[5] ));
    CCU2D add_7184_9 (.A0(\BUS_ADDR_INTERNAL[8]_adj_26 ), .B0(\BUS_ADDR_INTERNAL[8] ), 
          .C0(\BUS_currGrantID[0] ), .D0(\BUS_currGrantID[1] ), .A1(\BUS_ADDR_INTERNAL[9] ), 
          .B1(\BUS_ADDR_INTERNAL[9]_adj_27 ), .C1(\BUS_currGrantID[1] ), 
          .D1(\BUS_currGrantID[0] ), .CIN(n10160), .COUT(n10161));
    defparam add_7184_9.INIT0 = 16'hf530;
    defparam add_7184_9.INIT1 = 16'hf530;
    defparam add_7184_9.INJECT1_0 = "NO";
    defparam add_7184_9.INJECT1_1 = "NO";
    FD1S3DX state__i2 (.D(n10870), .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), 
            .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam state__i2.GSR = "DISABLED";
    PFUMX mux_472_i5 (.BLUT(Sprite_readData[4]), .ALUT(\otherData[4] ), 
          .C0(n11093), .Z(\BUS_DATA_INTERNAL[4] ));
    CCU2D add_7184_7 (.A0(\BUS_ADDR_INTERNAL[6]_adj_28 ), .B0(\BUS_ADDR_INTERNAL[6] ), 
          .C0(\BUS_currGrantID[0] ), .D0(\BUS_currGrantID[1] ), .A1(\BUS_ADDR_INTERNAL[7]_adj_29 ), 
          .B1(\BUS_ADDR_INTERNAL[7] ), .C1(\BUS_currGrantID[0] ), .D1(\BUS_currGrantID[1] ), 
          .CIN(n10159), .COUT(n10160));
    defparam add_7184_7.INIT0 = 16'hf530;
    defparam add_7184_7.INIT1 = 16'hf530;
    defparam add_7184_7.INJECT1_0 = "NO";
    defparam add_7184_7.INJECT1_1 = "NO";
    PFUMX mux_472_i4 (.BLUT(otherData[3]), .ALUT(n2372[3]), .C0(n1627), 
          .Z(\BUS_DATA_INTERNAL[3] ));
    FD1S3DX state__i1 (.D(n10540), .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam state__i1.GSR = "DISABLED";
    FD1S3AX yOffset_i7 (.D(yOffset_pre[7]), .CK(offsetLatchClockOrd), .Q(yOffset[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i7.GSR = "DISABLED";
    FD1S3AX yOffset_i6 (.D(yOffset_pre[6]), .CK(offsetLatchClockOrd), .Q(yOffset[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i6.GSR = "DISABLED";
    FD1S3AX yOffset_i5 (.D(yOffset_pre[5]), .CK(offsetLatchClockOrd), .Q(yOffset[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i5.GSR = "DISABLED";
    FD1S3AX yOffset_i4 (.D(yOffset_pre[4]), .CK(offsetLatchClockOrd), .Q(yOffset[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i4.GSR = "DISABLED";
    FD1S3AX yOffset_i3 (.D(yOffset_pre[3]), .CK(offsetLatchClockOrd), .Q(yOffset[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i3.GSR = "DISABLED";
    DPR16X4C n30442 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3032[0]), .DO1(n3032[1]));
    defparam n30442.initval = "0x0000000000000000";
    DPR16X4C n30402 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(VRAM_DATA[0]), .DO1(VRAM_DATA[1]));
    defparam n30402.initval = "0x0000000000000000";
    SPR16X4C Sprite_options15 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3383), .DO0(n3365), 
            .DO1(n3366), .DO2(n3367), .DO3(n3368));
    defparam Sprite_options15.initval = "0x0000000000000000";
    DPR16X4C n30422 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3029[0]), .DO1(n3029[1]));
    defparam n30422.initval = "0x0000000000000000";
    SPR16X4C Sprite_options14 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3383), .DO0(n3369), 
            .DO1(n3370), .DO2(n3371), .DO3(n3372));
    defparam Sprite_options14.initval = "0x0000000000000000";
    DPR16X4C n30462 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3035[0]), .DO1(n3035[1]));
    defparam n30462.initval = "0x0000000000000000";
    SPR16X4C Sprite_options13 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3383), .DO0(n3373), 
            .DO1(n3374), .DO2(n3375), .DO3(n3376));
    defparam Sprite_options13.initval = "0x0000000000000000";
    DPR16X4C n30400 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(VRAM_DATA[6]), .DO1(VRAM_DATA[7]), .DO2(VRAM_DATA[8]), 
            .DO3(VRAM_DATA[9]));
    defparam n30400.initval = "0x0000000000000000";
    SPR16X4C Sprite_options12 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3348), .DO0(n3330), 
            .DO1(n3331), .DO2(n3332), .DO3(n3333));
    defparam Sprite_options12.initval = "0x0000000000000000";
    DPR16X4C n30420 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3029[6]), .DO1(n3029[7]), .DO2(n3029[8]), .DO3(n3029[9]));
    defparam n30420.initval = "0x0000000000000000";
    SPR16X4C Sprite_options11 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3348), .DO0(n3334), 
            .DO1(n3335), .DO2(n3336), .DO3(n3337));
    defparam Sprite_options11.initval = "0x0000000000000000";
    DPR16X4C n30440 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3032[6]), .DO1(n3032[7]), .DO2(n3032[8]), .DO3(n3032[9]));
    defparam n30440.initval = "0x0000000000000000";
    SPR16X4C Sprite_options10 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3348), .DO0(n3338), 
            .DO1(n3339), .DO2(n3340), .DO3(n3341));
    defparam Sprite_options10.initval = "0x0000000000000000";
    DPR16X4C n30460 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(GND_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3035[6]), .DO1(n3035[7]), .DO2(n3035[8]), .DO3(n3035[9]));
    defparam n30460.initval = "0x0000000000000000";
    SPR16X4C Sprite_options9 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3382), .DO0(n3349), 
            .DO1(n3350), .DO2(n3351), .DO3(n3352));
    defparam Sprite_options9.initval = "0x0000000000000000";
    DPR16X4C n3039_d00 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3027[6]), .DO1(n3027[7]), .DO2(n3027[8]), .DO3(n3027[9]));
    defparam n3039_d00.initval = "0x0000000000000000";
    SPR16X4C Sprite_options8 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3382), .DO0(n3353), 
            .DO1(n3354), .DO2(n3355), .DO3(n3356));
    defparam Sprite_options8.initval = "0x0000000000000000";
    DPR16X4C n3040_d10 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3296), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3028[6]), .DO1(n3028[7]), .DO2(n3028[8]), .DO3(n3028[9]));
    defparam n3040_d10.initval = "0x0000000000000000";
    SPR16X4C Sprite_options7 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3382), .DO0(n3357), 
            .DO1(n3358), .DO2(n3359), .DO3(n3360));
    defparam Sprite_options7.initval = "0x0000000000000000";
    DPR16X4C n3041_d20 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3030[6]), .DO1(n3030[7]), .DO2(n3030[8]), .DO3(n3030[9]));
    defparam n3041_d20.initval = "0x0000000000000000";
    SPR16X4C Sprite_options6 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3347), .DO0(n3314), 
            .DO1(n3315), .DO2(n3316), .DO3(n3317));
    defparam Sprite_options6.initval = "0x0000000000000000";
    DPR16X4C n3042_d30 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3291), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3031[6]), .DO1(n3031[7]), .DO2(n3031[8]), .DO3(n3031[9]));
    defparam n3042_d30.initval = "0x0000000000000000";
    SPR16X4C Sprite_options5 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3347), .DO0(n3318), 
            .DO1(n3319), .DO2(n3320), .DO3(n3321));
    defparam Sprite_options5.initval = "0x0000000000000000";
    DPR16X4C n3043_d40 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3033[6]), .DO1(n3033[7]), .DO2(n3033[8]), .DO3(n3033[9]));
    defparam n3043_d40.initval = "0x0000000000000000";
    PFUMX mux_472_i3 (.BLUT(otherData[2]), .ALUT(n2372[2]), .C0(n1627), 
          .Z(\BUS_DATA_INTERNAL[2] ));
    CCU2D xPre_7__I_0_8 (.A0(xPre[6]), .B0(xOffset[6]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[7]), .B1(xOffset[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9979), .S0(x[6]), .S1(x[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(164[25:39])
    defparam xPre_7__I_0_8.INIT0 = 16'h5666;
    defparam xPre_7__I_0_8.INIT1 = 16'h5666;
    defparam xPre_7__I_0_8.INJECT1_0 = "NO";
    defparam xPre_7__I_0_8.INJECT1_1 = "NO";
    SPR16X4C Sprite_options0 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3382), .DO0(n3361), 
            .DO1(n3362), .DO2(n3363), .DO3(n3364));
    defparam Sprite_options0.initval = "0x0000000000000000";
    PFUMX mux_472_i2 (.BLUT(otherData[1]), .ALUT(n2372[1]), .C0(n1627), 
          .Z(\BUS_DATA_INTERNAL[1] ));
    DPR16X4C n3046_d70 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3037[6]), .DO1(n3037[7]), .DO2(n3037[8]), .DO3(n3037[9]));
    defparam n3046_d70.initval = "0x0000000000000000";
    CCU2D add_7184_5 (.A0(\BUS_ADDR_INTERNAL[4] ), .B0(\BUS_ADDR_INTERNAL[4]_adj_30 ), 
          .C0(\BUS_currGrantID[1] ), .D0(\BUS_currGrantID[0] ), .A1(\BUS_ADDR_INTERNAL[5] ), 
          .B1(\BUS_ADDR_INTERNAL[5]_adj_31 ), .C1(\BUS_currGrantID[1] ), 
          .D1(\BUS_currGrantID[0] ), .CIN(n10158), .COUT(n10159));
    defparam add_7184_5.INIT0 = 16'hf530;
    defparam add_7184_5.INIT1 = 16'hf530;
    defparam add_7184_5.INJECT1_0 = "NO";
    defparam add_7184_5.INJECT1_1 = "NO";
    FD1S3AX yOffset_i2 (.D(yOffset_pre[2]), .CK(offsetLatchClockOrd), .Q(yOffset[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i2.GSR = "DISABLED";
    DPR16X4C n3045_d60 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3306), 
            .RAD0(VCC_net), .RAD1(GND_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3036[6]), .DO1(n3036[7]), .DO2(n3036[8]), .DO3(n3036[9]));
    defparam n3045_d60.initval = "0x0000000000000000";
    SPR16X4C Sprite_options3 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3347), .DO0(n3326), 
            .DO1(n3327), .DO2(n3328), .DO3(n3329));
    defparam Sprite_options3.initval = "0x0000000000000000";
    SPR16X4C Sprite_options1 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3348), .DO0(n3342), 
            .DO1(n3343), .DO2(n3344), .DO3(n3345));
    defparam Sprite_options1.initval = "0x0000000000000000";
    CCU2D add_7184_3 (.A0(\BUS_ADDR_INTERNAL[2]_adj_32 ), .B0(\BUS_ADDR_INTERNAL[2] ), 
          .C0(\BUS_currGrantID[1] ), .D0(\BUS_currGrantID[0] ), .A1(\BUS_ADDR_INTERNAL[3]_adj_33 ), 
          .B1(\BUS_ADDR_INTERNAL[3] ), .C1(\BUS_currGrantID[0] ), .D1(\BUS_currGrantID[1] ), 
          .CIN(n10157), .COUT(n10158));
    defparam add_7184_3.INIT0 = 16'hf350;
    defparam add_7184_3.INIT1 = 16'hf530;
    defparam add_7184_3.INJECT1_0 = "NO";
    defparam add_7184_3.INJECT1_1 = "NO";
    SPR16X4C Sprite_options2 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3383), .DO0(n3377), 
            .DO1(n3378), .DO2(n3379), .DO3(n3380));
    defparam Sprite_options2.initval = "0x0000000000000000";
    DPR16X4C n3044_d50 (.DI0(GR_RE_DOUT[6]), .DI1(GR_RE_DOUT[7]), .DI2(GR_RE_DOUT[8]), 
            .DI3(GR_RE_DOUT[9]), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3034[6]), .DO1(n3034[7]), .DO2(n3034[8]), .DO3(n3034[9]));
    defparam n3044_d50.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes15 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3278), .DO0(n3260), 
            .DO1(n3261), .DO2(n3262), .DO3(n3263));
    defparam Sprite_sizes15.initval = "0x0000000000000000";
    CCU2D xPre_7__I_0_6 (.A0(xPre[4]), .B0(xOffset[4]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[5]), .B1(xOffset[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9978), .COUT(n9979), .S0(x[4]), .S1(x[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(164[25:39])
    defparam xPre_7__I_0_6.INIT0 = 16'h5666;
    defparam xPre_7__I_0_6.INIT1 = 16'h5666;
    defparam xPre_7__I_0_6.INJECT1_0 = "NO";
    defparam xPre_7__I_0_6.INJECT1_1 = "NO";
    CCU2D add_7184_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n12277), .B1(n12344), .C1(n12292), .D1(GND_net), .COUT(n10157));
    defparam add_7184_1.INIT0 = 16'hF000;
    defparam add_7184_1.INIT1 = 16'hb848;
    defparam add_7184_1.INJECT1_0 = "NO";
    defparam add_7184_1.INJECT1_1 = "NO";
    PFUMX mux_472_i1 (.BLUT(otherData[0]), .ALUT(n2372[0]), .C0(n1627), 
          .Z(\BUS_DATA_INTERNAL[0] ));
    SPR16X4C Sprite_sizes14 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3278), .DO0(n3264), 
            .DO1(n3265), .DO2(n3266), .DO3(n3267));
    defparam Sprite_sizes14.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes13 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3278), .DO0(n3268), 
            .DO1(n3269), .DO2(n3270), .DO3(n3271));
    defparam Sprite_sizes13.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes12 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3243), .DO0(n3225), 
            .DO1(n3226), .DO2(n3227), .DO3(n3228));
    defparam Sprite_sizes12.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes11 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3243), .DO0(n3229), 
            .DO1(n3230), .DO2(n3231), .DO3(n3232));
    defparam Sprite_sizes11.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes10 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3243), .DO0(n3233), 
            .DO1(n3234), .DO2(n3235), .DO3(n3236));
    defparam Sprite_sizes10.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes9 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3277), .DO0(n3244), 
            .DO1(n3245), .DO2(n3246), .DO3(n3247));
    defparam Sprite_sizes9.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes8 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3277), .DO0(n3248), 
            .DO1(n3249), .DO2(n3250), .DO3(n3251));
    defparam Sprite_sizes8.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes7 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3277), .DO0(n3252), 
            .DO1(n3253), .DO2(n3254), .DO3(n3255));
    defparam Sprite_sizes7.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes6 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3242), .DO0(n3209), 
            .DO1(n3210), .DO2(n3211), .DO3(n3212));
    defparam Sprite_sizes6.initval = "0x0000000000000000";
    L6MUX21 i8257 (.D0(n11147), .D1(n11148), .SD(n12269), .Z(n11149));
    SPR16X4C Sprite_sizes5 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3242), .DO0(n3213), 
            .DO1(n3214), .DO2(n3215), .DO3(n3216));
    defparam Sprite_sizes5.initval = "0x0000000000000000";
    L6MUX21 i8264 (.D0(n11154), .D1(n11155), .SD(n12269), .Z(n11156));
    L6MUX21 i8208 (.D0(n11098), .D1(n11099), .SD(n12269), .Z(n11100));
    LUT4 currColor_1__bdd_3_lut (.A(currColor[1]), .B(currColor[2]), .C(currColor[0]), 
         .Z(n12049)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;
    defparam currColor_1__bdd_3_lut.init = 16'h6c6c;
    SPR16X4C Sprite_sizes0 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3277), .DO0(n3256), 
            .DO1(n3257), .DO2(n3258), .DO3(n3259));
    defparam Sprite_sizes0.initval = "0x0000000000000000";
    L6MUX21 i8271 (.D0(n11161), .D1(n11162), .SD(n12269), .Z(n11163));
    L6MUX21 i8278 (.D0(n11168), .D1(n11169), .SD(n12269), .Z(n11170));
    SPR16X4C Sprite_sizes3 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3242), .DO0(n3221), 
            .DO1(n3222), .DO2(n3223), .DO3(n3224));
    defparam Sprite_sizes3.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes1 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3243), .DO0(n3237), 
            .DO1(n3238), .DO2(n3239), .DO3(n3240));
    defparam Sprite_sizes1.initval = "0x0000000000000000";
    SPR16X4C Sprite_sizes2 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), .DI2(BUS_data[14]), 
            .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3278), .DO0(n3272), 
            .DO1(n3273), .DO2(n3274), .DO3(n3275));
    defparam Sprite_sizes2.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions15 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3173), .DO0(n3155), 
            .DO1(n3156), .DO2(n3157), .DO3(n3158));
    defparam Sprite_positions15.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions14 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3173), .DO0(n3159), 
            .DO1(n3160), .DO2(n3161), .DO3(n3162));
    defparam Sprite_positions14.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions13 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3173), .DO0(n3163), 
            .DO1(n3164), .DO2(n3165), .DO3(n3166));
    defparam Sprite_positions13.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions12 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3138), .DO0(n3120), 
            .DO1(n3121), .DO2(n3122), .DO3(n3123));
    defparam Sprite_positions12.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions11 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3138), .DO0(n3124), 
            .DO1(n3125), .DO2(n3126), .DO3(n3127));
    defparam Sprite_positions11.initval = "0x0000000000000000";
    L6MUX21 i8215 (.D0(n11105), .D1(n11106), .SD(n12269), .Z(n11107));
    SPR16X4C Sprite_positions10 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3138), .DO0(n3128), 
            .DO1(n3129), .DO2(n3130), .DO3(n3131));
    defparam Sprite_positions10.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions9 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3172), .DO0(n3139), 
            .DO1(n3140), .DO2(n3141), .DO3(n3142));
    defparam Sprite_positions9.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions8 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3172), .DO0(n3143), 
            .DO1(n3144), .DO2(n3145), .DO3(n3146));
    defparam Sprite_positions8.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions7 (.DI0(BUS_data[8]), .DI1(BUS_data[9]), .DI2(BUS_data[10]), 
            .DI3(BUS_data[11]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3172), .DO0(n3147), 
            .DO1(n3148), .DO2(n3149), .DO3(n3150));
    defparam Sprite_positions7.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions6 (.DI0(BUS_data[0]), .DI1(BUS_data[1]), .DI2(BUS_data[2]), 
            .DI3(BUS_data[3]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3137), .DO0(n3104), 
            .DO1(n3105), .DO2(n3106), .DO3(n3107));
    defparam Sprite_positions6.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions5 (.DI0(BUS_data[4]), .DI1(BUS_data[5]), .DI2(BUS_data[6]), 
            .DI3(BUS_data[7]), .AD0(n12253), .AD1(n12264), .AD2(n12259), 
            .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3137), .DO0(n3108), 
            .DO1(n3109), .DO2(n3110), .DO3(n3111));
    defparam Sprite_positions5.initval = "0x0000000000000000";
    L6MUX21 i8300 (.D0(n11190), .D1(n11191), .SD(n12269), .Z(n11192));
    CCU2D add_7186_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10136), 
          .S0(n2129));
    defparam add_7186_cout.INIT0 = 16'h0000;
    defparam add_7186_cout.INIT1 = 16'h0000;
    defparam add_7186_cout.INJECT1_0 = "NO";
    defparam add_7186_cout.INJECT1_1 = "NO";
    DPR16X4C n3044_d52 (.DI0(GR_RE_DOUT[0]), .DI1(GR_RE_DOUT[1]), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(currColor_lat[0]), .WAD1(currColor_lat[1]), 
            .WAD2(GND_net), .WAD3(GND_net), .WCK(LOGIC_CLOCK), .WRE(n3301), 
            .RAD0(GND_net), .RAD1(VCC_net), .RAD2(GND_net), .RAD3(GND_net), 
            .DO0(n3034[0]), .DO1(n3034[1]));
    defparam n3044_d52.initval = "0x0000000000000000";
    SPR16X4C Sprite_positions0 (.DI0(BUS_data[12]), .DI1(BUS_data[13]), 
            .DI2(BUS_data[14]), .DI3(BUS_data[15]), .AD0(n12253), .AD1(n12264), 
            .AD2(n12259), .AD3(n12247), .CK(LOGIC_CLOCK), .WRE(n3172), 
            .DO0(n3151), .DO1(n3152), .DO2(n3153), .DO3(n3154));
    defparam Sprite_positions0.initval = "0x0000000000000000";
    L6MUX21 i8313 (.D0(n11203), .D1(n11204), .SD(n12269), .Z(n11205));
    FD1P3AX currValue_i0_i0 (.D(BUS_data[0]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i0.GSR = "DISABLED";
    FD1P3DX currColor_683__i0 (.D(n27[0]), .SP(LOGIC_CLOCK_enable_178), 
            .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), .Q(currColor[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_683__i0.GSR = "DISABLED";
    FD1S3AX yOffset_i1 (.D(yOffset_pre[1]), .CK(offsetLatchClockOrd), .Q(yOffset[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam yOffset_i1.GSR = "DISABLED";
    CCU2D add_7186_13 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n10135), .COUT(n10136));
    defparam add_7186_13.INIT0 = 16'heeee;
    defparam add_7186_13.INIT1 = 16'heeee;
    defparam add_7186_13.INJECT1_0 = "NO";
    defparam add_7186_13.INJECT1_1 = "NO";
    L6MUX21 i8329 (.D0(n11219), .D1(n11220), .SD(n12269), .Z(n11221));
    CCU2D add_7186_11 (.A0(n13158), .B0(n12344), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), 
          .D1(n12309), .CIN(n10134), .COUT(n10135));
    defparam add_7186_11.INIT0 = 16'h8888;
    defparam add_7186_11.INIT1 = 16'hff20;
    defparam add_7186_11.INJECT1_0 = "NO";
    defparam add_7186_11.INJECT1_1 = "NO";
    CCU2D add_7186_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n13150), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16]_adj_19 ), 
          .D1(n13151), .CIN(n10133), .COUT(n10134));
    defparam add_7186_9.INIT0 = 16'hff51;
    defparam add_7186_9.INIT1 = 16'hff51;
    defparam add_7186_9.INJECT1_0 = "NO";
    defparam add_7186_9.INJECT1_1 = "NO";
    FD1P3AX reset_344 (.D(reset_N_670), .SP(state_7__N_322), .CK(LOGIC_CLOCK), 
            .Q(reset)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam reset_344.GSR = "DISABLED";
    L6MUX21 i8222 (.D0(n11112), .D1(n11113), .SD(n12269), .Z(n11114));
    CCU2D add_7186_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n13155), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n13157), 
          .CIN(n10132), .COUT(n10133));
    defparam add_7186_7.INIT0 = 16'h00ae;
    defparam add_7186_7.INIT1 = 16'h00ae;
    defparam add_7186_7.INJECT1_0 = "NO";
    defparam add_7186_7.INJECT1_1 = "NO";
    CCU2D add_7186_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n13156), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n13142), 
          .CIN(n10131), .COUT(n10132));
    defparam add_7186_5.INIT0 = 16'h00ae;
    defparam add_7186_5.INIT1 = 16'h00ae;
    defparam add_7186_5.INJECT1_0 = "NO";
    defparam add_7186_5.INJECT1_1 = "NO";
    CCU2D add_7186_3 (.A0(\BUS_ADDR_INTERNAL[9] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13144), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n13143), 
          .CIN(n10130), .COUT(n10131));
    defparam add_7186_3.INIT0 = 16'h00dc;
    defparam add_7186_3.INIT1 = 16'h00ae;
    defparam add_7186_3.INJECT1_0 = "NO";
    defparam add_7186_3.INJECT1_1 = "NO";
    CCU2D add_7186_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), 
          .D1(n13154), .COUT(n10130));
    defparam add_7186_1.INIT0 = 16'hF000;
    defparam add_7186_1.INIT1 = 16'h00ae;
    defparam add_7186_1.INJECT1_0 = "NO";
    defparam add_7186_1.INJECT1_1 = "NO";
    FD1P3DX latchForce_365 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_49), 
            .CK(LOGIC_CLOCK), .CD(n12219), .Q(latchForce)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam latchForce_365.GSR = "DISABLED";
    L6MUX21 i8229 (.D0(n11119), .D1(n11120), .SD(n12269), .Z(n11121));
    L6MUX21 i8236 (.D0(n11126), .D1(n11127), .SD(n12269), .Z(n11128));
    L6MUX21 i8243 (.D0(n11133), .D1(n11134), .SD(n12269), .Z(n11135));
    L6MUX21 i8438 (.D0(n11328), .D1(n11329), .SD(n12269), .Z(n11330));
    L6MUX21 i8445 (.D0(n11335), .D1(n11336), .SD(n12269), .Z(n11337));
    FD1P3AX xOffset_pre_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i7.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i6.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i5.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i4.GSR = "DISABLED";
    L6MUX21 i8250 (.D0(n11140), .D1(n11141), .SD(n12269), .Z(n11142));
    PFUMX i8206 (.BLUT(n11094), .ALUT(n11095), .C0(n12263), .Z(n11098));
    FD1P3AX xOffset_pre_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i3.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i2.GSR = "DISABLED";
    FD1P3AX xOffset_pre_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_71), 
            .CK(LOGIC_CLOCK), .Q(xOffset_pre[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam xOffset_pre_i0_i1.GSR = "DISABLED";
    PFUMX i8207 (.BLUT(n11096), .ALUT(n11097), .C0(n12263), .Z(n11099));
    PFUMX i8262 (.BLUT(n11150), .ALUT(n11151), .C0(n12263), .Z(n11154));
    PFUMX i8263 (.BLUT(n11152), .ALUT(n11153), .C0(n12263), .Z(n11155));
    PFUMX i8269 (.BLUT(n11157), .ALUT(n11158), .C0(n12263), .Z(n11161));
    PFUMX i8270 (.BLUT(n11159), .ALUT(n11160), .C0(n12263), .Z(n11162));
    PFUMX i8276 (.BLUT(n11164), .ALUT(n11165), .C0(n12263), .Z(n11168));
    PFUMX i8277 (.BLUT(n11166), .ALUT(n11167), .C0(n12263), .Z(n11169));
    CCU2D add_7188_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10084), .S1(n1921));
    defparam add_7188_21.INIT0 = 16'heeee;
    defparam add_7188_21.INIT1 = 16'h0000;
    defparam add_7188_21.INJECT1_0 = "NO";
    defparam add_7188_21.INJECT1_1 = "NO";
    CCU2D xPre_7__I_0_4 (.A0(xPre[2]), .B0(xOffset[2]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[3]), .B1(xOffset[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9977), .COUT(n9978), .S0(x[2]), .S1(x[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(164[25:39])
    defparam xPre_7__I_0_4.INIT0 = 16'h5666;
    defparam xPre_7__I_0_4.INIT1 = 16'h5666;
    defparam xPre_7__I_0_4.INJECT1_0 = "NO";
    defparam xPre_7__I_0_4.INJECT1_1 = "NO";
    PFUMX i8281 (.BLUT(n11171), .ALUT(n11172), .C0(n12263), .Z(Sprite_readData_15__N_417[14]));
    FD1P3AX yOffset_pre_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i1.GSR = "DISABLED";
    CCU2D add_7188_19 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[18] ), .D0(n12309), .A1(\BUS_currGrantID[0] ), 
          .B1(\BUS_currGrantID[1] ), .C1(GND_net), .D1(GND_net), .CIN(n10083), 
          .COUT(n10084));
    defparam add_7188_19.INIT0 = 16'hff20;
    defparam add_7188_19.INIT1 = 16'heeee;
    defparam add_7188_19.INJECT1_0 = "NO";
    defparam add_7188_19.INJECT1_1 = "NO";
    PFUMX i8284 (.BLUT(n11174), .ALUT(n11175), .C0(n12263), .Z(Sprite_readData_15__N_417[15]));
    CCU2D add_7188_17 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[16]_adj_19 ), .D0(n13151), .A1(n13158), 
          .B1(n12344), .C1(GND_net), .D1(GND_net), .CIN(n10082), .COUT(n10083));
    defparam add_7188_17.INIT0 = 16'h00ae;
    defparam add_7188_17.INIT1 = 16'h8888;
    defparam add_7188_17.INJECT1_0 = "NO";
    defparam add_7188_17.INJECT1_1 = "NO";
    PFUMX i8287 (.BLUT(n11177), .ALUT(n11178), .C0(n12263), .Z(Sprite_readData_15__N_417[0]));
    CCU2D add_7188_15 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[14] ), .D0(n13157), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[15] ), .D1(n13150), 
          .CIN(n10081), .COUT(n10082));
    defparam add_7188_15.INIT0 = 16'h00ae;
    defparam add_7188_15.INIT1 = 16'h00ae;
    defparam add_7188_15.INJECT1_0 = "NO";
    defparam add_7188_15.INJECT1_1 = "NO";
    CCU2D add_7188_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[12] ), .D0(n13142), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[13] ), .D1(n13155), 
          .CIN(n10080), .COUT(n10081));
    defparam add_7188_13.INIT0 = 16'h00ae;
    defparam add_7188_13.INIT1 = 16'h00ae;
    defparam add_7188_13.INJECT1_0 = "NO";
    defparam add_7188_13.INJECT1_1 = "NO";
    PFUMX i8290 (.BLUT(n11180), .ALUT(n11181), .C0(n12263), .Z(Sprite_readData_15__N_417[1]));
    CCU2D add_7188_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[10] ), .D0(n13143), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[11] ), .D1(n13156), 
          .CIN(n10079), .COUT(n10080));
    defparam add_7188_11.INIT0 = 16'hff51;
    defparam add_7188_11.INIT1 = 16'h00ae;
    defparam add_7188_11.INJECT1_0 = "NO";
    defparam add_7188_11.INJECT1_1 = "NO";
    CCU2D add_1231_9 (.A0(x[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n9995), 
          .S0(currAddress_17__N_506[8]), .S1(currAddress_17__N_506[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[150:167])
    defparam add_1231_9.INIT0 = 16'h5aaa;
    defparam add_1231_9.INIT1 = 16'h0000;
    defparam add_1231_9.INJECT1_0 = "NO";
    defparam add_1231_9.INJECT1_1 = "NO";
    CCU2D add_7188_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[8] ), .D0(n13154), .A1(\BUS_ADDR_INTERNAL[9] ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13144), 
          .CIN(n10078), .COUT(n10079));
    defparam add_7188_9.INIT0 = 16'h00ae;
    defparam add_7188_9.INIT1 = 16'h00dc;
    defparam add_7188_9.INJECT1_0 = "NO";
    defparam add_7188_9.INJECT1_1 = "NO";
    FD1P3AX yOffset_pre_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i2.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i3.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i4.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i5.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i6.GSR = "DISABLED";
    FD1P3AX yOffset_pre_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_78), 
            .CK(LOGIC_CLOCK), .Q(yOffset_pre[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam yOffset_pre_i0_i7.GSR = "DISABLED";
    FD1P3AX latchMode_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_81), 
            .CK(LOGIC_CLOCK), .Q(latchMode[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam latchMode_i0_i1.GSR = "DISABLED";
    CCU2D add_1231_7 (.A0(x[5]), .B0(x[6]), .C0(GND_net), .D0(GND_net), 
          .A1(x[6]), .B1(x[7]), .C1(GND_net), .D1(GND_net), .CIN(n9994), 
          .COUT(n9995), .S0(currAddress_17__N_506[6]), .S1(currAddress_17__N_506[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[150:167])
    defparam add_1231_7.INIT0 = 16'h5666;
    defparam add_1231_7.INIT1 = 16'h5666;
    defparam add_1231_7.INJECT1_0 = "NO";
    defparam add_1231_7.INJECT1_1 = "NO";
    PFUMX i8293 (.BLUT(n11183), .ALUT(n11184), .C0(n12263), .Z(Sprite_readData_15__N_417[2]));
    CCU2D add_7188_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[6] ), .D0(n13146), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[7] ), .D1(n13147), 
          .CIN(n10077), .COUT(n10078));
    defparam add_7188_7.INIT0 = 16'h00ae;
    defparam add_7188_7.INIT1 = 16'h00ae;
    defparam add_7188_7.INJECT1_0 = "NO";
    defparam add_7188_7.INJECT1_1 = "NO";
    FD1P3AX latchMode_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_81), 
            .CK(LOGIC_CLOCK), .Q(latchMode[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam latchMode_i0_i2.GSR = "DISABLED";
    FD1P3AX latchMode_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_81), 
            .CK(LOGIC_CLOCK), .Q(latchMode[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam latchMode_i0_i3.GSR = "DISABLED";
    FD1S3AX xOffset_i1 (.D(xOffset_pre[1]), .CK(offsetLatchClockOrd), .Q(xOffset[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i1.GSR = "DISABLED";
    CCU2D add_7188_5 (.A0(\BUS_ADDR_INTERNAL[4] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13153), .A1(\BUS_ADDR_INTERNAL[5] ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13145), 
          .CIN(n10076), .COUT(n10077));
    defparam add_7188_5.INIT0 = 16'h00dc;
    defparam add_7188_5.INIT1 = 16'h00dc;
    defparam add_7188_5.INJECT1_0 = "NO";
    defparam add_7188_5.INJECT1_1 = "NO";
    CCU2D add_7188_3 (.A0(\BUS_ADDR_INTERNAL[2] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13152), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[3] ), .D1(n13148), 
          .CIN(n10075), .COUT(n10076));
    defparam add_7188_3.INIT0 = 16'h00dc;
    defparam add_7188_3.INIT1 = 16'h00ae;
    defparam add_7188_3.INJECT1_0 = "NO";
    defparam add_7188_3.INJECT1_1 = "NO";
    FD1S3AX xOffset_i2 (.D(xOffset_pre[2]), .CK(offsetLatchClockOrd), .Q(xOffset[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i2.GSR = "DISABLED";
    FD1S3AX xOffset_i3 (.D(xOffset_pre[3]), .CK(offsetLatchClockOrd), .Q(xOffset[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i3.GSR = "DISABLED";
    FD1S3AX xOffset_i4 (.D(xOffset_pre[4]), .CK(offsetLatchClockOrd), .Q(xOffset[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i4.GSR = "DISABLED";
    FD1S3AX xOffset_i5 (.D(xOffset_pre[5]), .CK(offsetLatchClockOrd), .Q(xOffset[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i5.GSR = "DISABLED";
    FD1S3AX xOffset_i6 (.D(xOffset_pre[6]), .CK(offsetLatchClockOrd), .Q(xOffset[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i6.GSR = "DISABLED";
    FD1S3AX xOffset_i7 (.D(xOffset_pre[7]), .CK(offsetLatchClockOrd), .Q(xOffset[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(176[3] 179[10])
    defparam xOffset_i7.GSR = "DISABLED";
    CCU2D add_1231_5 (.A0(x[3]), .B0(x[4]), .C0(GND_net), .D0(GND_net), 
          .A1(x[4]), .B1(x[5]), .C1(GND_net), .D1(GND_net), .CIN(n9993), 
          .COUT(n9994), .S0(currAddress_17__N_506[4]), .S1(currAddress_17__N_506[5]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[150:167])
    defparam add_1231_5.INIT0 = 16'h5666;
    defparam add_1231_5.INIT1 = 16'h5666;
    defparam add_1231_5.INJECT1_0 = "NO";
    defparam add_1231_5.INJECT1_1 = "NO";
    PFUMX i8213 (.BLUT(n11101), .ALUT(n11102), .C0(n12263), .Z(n11105));
    CCU2D add_7188_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n12292), .B1(n12344), .C1(n13139), .D1(n12299), .COUT(n10075));
    defparam add_7188_1.INIT0 = 16'hF000;
    defparam add_7188_1.INIT1 = 16'h4448;
    defparam add_7188_1.INJECT1_0 = "NO";
    defparam add_7188_1.INJECT1_1 = "NO";
    CCU2D add_1231_3 (.A0(x[1]), .B0(x[2]), .C0(GND_net), .D0(GND_net), 
          .A1(x[2]), .B1(x[3]), .C1(GND_net), .D1(GND_net), .CIN(n9992), 
          .COUT(n9993), .S0(currAddress_17__N_506[2]), .S1(currAddress_17__N_506[3]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[150:167])
    defparam add_1231_3.INIT0 = 16'h5666;
    defparam add_1231_3.INIT1 = 16'h5666;
    defparam add_1231_3.INJECT1_0 = "NO";
    defparam add_1231_3.INJECT1_1 = "NO";
    PFUMX i8214 (.BLUT(n11103), .ALUT(n11104), .C0(n12263), .Z(n11106));
    LUT4 i1_4_lut (.A(n10309), .B(n11156), .C(Sprite_readData_15__N_417[13]), 
         .D(n12265), .Z(\MDM_data[13] )) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h5044;
    CCU2D add_1231_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[0]), .B1(xOffset[0]), .C1(x[1]), .D1(GND_net), .COUT(n9992), 
          .S1(currAddress_17__N_506[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[150:167])
    defparam add_1231_1.INIT0 = 16'hF000;
    defparam add_1231_1.INIT1 = 16'h9696;
    defparam add_1231_1.INJECT1_0 = "NO";
    defparam add_1231_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_150 (.A(n10309), .B(n11163), .C(Sprite_readData_15__N_417[14]), 
         .D(n12265), .Z(\MDM_data[14] )) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    defparam i1_4_lut_adj_150.init = 16'h5044;
    LUT4 i2_4_lut (.A(n13), .B(n12261), .C(n100), .D(\BUS_DATA_INTERNAL[15] ), 
         .Z(BUS_data[15])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    defparam i2_4_lut.init = 16'hfefa;
    LUT4 i1_2_lut_4_lut (.A(n12292), .B(n12269), .C(n12218), .D(n4537), 
         .Z(n3138)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_4_lut (.A(state[0]), .B(BUS_DONE), .C(state[1]), .D(n12331), 
         .Z(n10540)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((D)+!C))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h0058;
    PFUMX i8298 (.BLUT(n11186), .ALUT(n11187), .C0(n12263), .Z(n11190));
    LUT4 i1_2_lut_4_lut_adj_151 (.A(n12292), .B(n12269), .C(n12218), .D(n4541), 
         .Z(n3173)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_151.init = 16'h0100;
    LUT4 i2_4_lut_adj_152 (.A(BUS_DONE_OUT_N_627), .B(n12230), .C(n63), 
         .D(n1184), .Z(n10846)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(323[4] 373[11])
    defparam i2_4_lut_adj_152.init = 16'hbfff;
    LUT4 BUS_VALID_N_480_I_0_2_lut (.A(BUS_VALID_N_480), .B(BUS_DONE_OUT_N_626), 
         .Z(BUS_DONE_OUT_N_627)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(352[11:65])
    defparam BUS_VALID_N_480_I_0_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_4_lut_adj_153 (.A(n12292), .B(n12269), .C(n12218), .D(n4545), 
         .Z(n3172)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_153.init = 16'h0100;
    LUT4 i4671_4_lut (.A(Sprite_readData[8]), .B(n3790), .C(GR_WR_DOUT[8]), 
         .D(n1956), .Z(\MDM_data[8] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(283[18:101])
    defparam i4671_4_lut.init = 16'h3022;
    PFUMX i8299 (.BLUT(n11188), .ALUT(n11189), .C0(n12263), .Z(n11191));
    LUT4 i4680_4_lut (.A(Sprite_readData[9]), .B(n3790), .C(GR_WR_DOUT[9]), 
         .D(n1956), .Z(\MDM_data[9] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(283[18:101])
    defparam i4680_4_lut.init = 16'h3022;
    PFUMX i8303 (.BLUT(n11193), .ALUT(n11194), .C0(n12263), .Z(Sprite_readData_15__N_417[3]));
    CCU2D xPre_7__I_0_2 (.A0(xPre[0]), .B0(xOffset[0]), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[1]), .B1(xOffset[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n9977), .S1(x[1]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(164[25:39])
    defparam xPre_7__I_0_2.INIT0 = 16'h7000;
    defparam xPre_7__I_0_2.INIT1 = 16'h5666;
    defparam xPre_7__I_0_2.INJECT1_0 = "NO";
    defparam xPre_7__I_0_2.INJECT1_1 = "NO";
    CCU2D add_1230_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10042), 
          .S0(currAddress_17__N_488[17]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[112:132])
    defparam add_1230_cout.INIT0 = 16'h0000;
    defparam add_1230_cout.INIT1 = 16'h0000;
    defparam add_1230_cout.INJECT1_0 = "NO";
    defparam add_1230_cout.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_154 (.A(n10309), .B(n11135), .C(Sprite_readData_15__N_417[10]), 
         .D(n12265), .Z(\MDM_data[10] )) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    defparam i1_4_lut_adj_154.init = 16'h5044;
    CCU2D add_1230_8 (.A0(y[7]), .B0(n4), .C0(n10348), .D0(GND_net), 
          .A1(y[7]), .B1(n4), .C1(GND_net), .D1(GND_net), .CIN(n10041), 
          .COUT(n10042), .S0(currAddress_17__N_488[15]), .S1(currAddress_17__N_488[16]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[112:132])
    defparam add_1230_8.INIT0 = 16'h9696;
    defparam add_1230_8.INIT1 = 16'h9666;
    defparam add_1230_8.INJECT1_0 = "NO";
    defparam add_1230_8.INJECT1_1 = "NO";
    LUT4 n12092_bdd_3_lut (.A(n12092), .B(VRAM_WC), .C(state[1]), .Z(VRAM_WC_N_598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n12092_bdd_3_lut.init = 16'hcaca;
    CCU2D add_1230_6 (.A0(y[5]), .B0(currRowOffset[0]), .C0(y[4]), .D0(GND_net), 
          .A1(currRowOffset[1]), .B1(n4_adj_1294), .C1(n162[5]), .D1(GND_net), 
          .CIN(n10040), .COUT(n10041), .S0(currAddress_17__N_488[13]), 
          .S1(currAddress_17__N_488[14]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[112:132])
    defparam add_1230_6.INIT0 = 16'h9696;
    defparam add_1230_6.INIT1 = 16'h9696;
    defparam add_1230_6.INJECT1_0 = "NO";
    defparam add_1230_6.INJECT1_1 = "NO";
    CCU2D yPre_7__I_0_7 (.A0(yOffset[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(yOffset[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9983), .COUT(n9984), .S0(y[5]), .S1(y[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(165[24:38])
    defparam yPre_7__I_0_7.INIT0 = 16'hfaaa;
    defparam yPre_7__I_0_7.INIT1 = 16'hfaaa;
    defparam yPre_7__I_0_7.INJECT1_0 = "NO";
    defparam yPre_7__I_0_7.INJECT1_1 = "NO";
    CCU2D add_1230_4 (.A0(y[2]), .B0(y[3]), .C0(GND_net), .D0(GND_net), 
          .A1(y[3]), .B1(y[4]), .C1(GND_net), .D1(GND_net), .CIN(n10039), 
          .COUT(n10040), .S0(currAddress_17__N_488[11]), .S1(currAddress_17__N_488[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[112:132])
    defparam add_1230_4.INIT0 = 16'h5666;
    defparam add_1230_4.INIT1 = 16'h5666;
    defparam add_1230_4.INJECT1_0 = "NO";
    defparam add_1230_4.INJECT1_1 = "NO";
    LUT4 i7326_4_lut_4_lut_rep_343 (.A(\BUS_currGrantID[1] ), .B(\BUS_currGrantID[0] ), 
         .C(\BUS_ADDR_INTERNAL[17] ), .D(BUS_ADDR_INTERNAL[17]), .Z(n13158)) /* synthesis lut_function=(A (B+!(C))+!A !(B (D))) */ ;
    defparam i7326_4_lut_4_lut_rep_343.init = 16'h9bdf;
    LUT4 i8729_2_lut_rep_303_3_lut_4_lut (.A(\BUS_currGrantID[1] ), .B(\BUS_currGrantID[0] ), 
         .C(\BUS_ADDR_INTERNAL[17] ), .D(BUS_ADDR_INTERNAL[17]), .Z(n12329)) /* synthesis lut_function=(!(A (B+!(C))+!A !((D)+!B))) */ ;
    defparam i8729_2_lut_rep_303_3_lut_4_lut.init = 16'h7531;
    CCU2D yPre_7__I_0_9 (.A0(yOffset[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n9984), .S0(y[7]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(165[24:38])
    defparam yPre_7__I_0_9.INIT0 = 16'hfaaa;
    defparam yPre_7__I_0_9.INIT1 = 16'h0000;
    defparam yPre_7__I_0_9.INJECT1_0 = "NO";
    defparam yPre_7__I_0_9.INJECT1_1 = "NO";
    FD1P3DX xPre_681__i1 (.D(n37[1]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[1])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i1.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_4_lut (.A(n12219), .B(n1184), .C(n12230), .D(n12226), 
         .Z(LOGIC_CLOCK_enable_78)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 i1_4_lut_adj_155 (.A(n10309), .B(n11142), .C(Sprite_readData_15__N_417[11]), 
         .D(n12265), .Z(\MDM_data[11] )) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    defparam i1_4_lut_adj_155.init = 16'h5044;
    LUT4 i1_2_lut_3_lut_3_lut (.A(n12219), .B(n1627), .C(n13141), .Z(n3790)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam i1_2_lut_3_lut_3_lut.init = 16'hfefe;
    LUT4 i4571_4_lut (.A(BUS_transferState[3]), .B(LOGIC_CLOCK_enable_26), 
         .C(n8), .D(n12228), .Z(LOGIC_CLOCK_enable_10)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(323[4] 373[11])
    defparam i4571_4_lut.init = 16'hdccc;
    LUT4 i3_3_lut_4_lut (.A(n12215), .B(n1956), .C(n12_adj_1295), .D(n1627), 
         .Z(n13)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0020;
    LUT4 state_2__bdd_4_lut (.A(state[2]), .B(state[4]), .C(VRAM_WC), 
         .D(state[0]), .Z(n12092)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C (D))+!B !((D)+!C))) */ ;
    defparam state_2__bdd_4_lut.init = 16'he0b2;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(n12219), .B(n1956), .C(n1627), 
         .D(n13141), .Z(n10309)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'hfffe;
    PFUMX i8306 (.BLUT(n11196), .ALUT(n11197), .C0(n12263), .Z(Sprite_readData_15__N_417[4]));
    LUT4 i1_2_lut_3_lut_4_lut (.A(n12224), .B(n12219), .C(n12244), .D(n12265), 
         .Z(n3347)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D add_1230_2 (.A0(currAddress_17__N_488[8]), .B0(y[1]), .C0(GND_net), 
          .D0(GND_net), .A1(y[1]), .B1(y[2]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10039), .S1(currAddress_17__N_488[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[112:132])
    defparam add_1230_2.INIT0 = 16'h7000;
    defparam add_1230_2.INIT1 = 16'h5666;
    defparam add_1230_2.INJECT1_0 = "NO";
    defparam add_1230_2.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_156 (.A(n12224), .B(n12219), .C(n4541), 
         .D(n12265), .Z(n3383)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_156.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_157 (.A(n12224), .B(n12219), .C(n4537), 
         .D(n12265), .Z(n3348)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_157.init = 16'h1000;
    LUT4 i9_4_lut (.A(n12332), .B(n18), .C(n12352), .D(n11052), .Z(n10898)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+(D))+!B))) */ ;
    defparam i9_4_lut.init = 16'h080c;
    LUT4 i1_2_lut_3_lut_4_lut_adj_158 (.A(n12224), .B(n12219), .C(n4545), 
         .D(n12265), .Z(n3382)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_158.init = 16'h1000;
    LUT4 BUS_DONE_OUT_N_625_bdd_4_lut (.A(n10846), .B(n13141), .C(LOGIC_CLOCK_enable_26), 
         .D(BUS_transferState[3]), .Z(n12157)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam BUS_DONE_OUT_N_625_bdd_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_2_lut_4_lut (.A(BUS_VALID_N_480), .B(n12222), .C(n2129), 
         .D(LOGIC_CLOCK_enable_49), .Z(LOGIC_CLOCK_enable_81)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (B+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam i1_2_lut_2_lut_4_lut.init = 16'h3b00;
    LUT4 i1_2_lut_rep_189_2_lut_4_lut (.A(BUS_VALID_N_480), .B(n12222), 
         .C(n2129), .D(n13141), .Z(n12215)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (B+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam i1_2_lut_rep_189_2_lut_4_lut.init = 16'h003b;
    LUT4 n12158_bdd_2_lut_rep_192_4_lut (.A(BUS_VALID_N_480), .B(n12222), 
         .C(n2129), .D(n12224), .Z(n12218)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam n12158_bdd_2_lut_rep_192_4_lut.init = 16'hffc4;
    LUT4 inv_38_i7_1_lut (.A(xPre[6]), .Z(n280[6])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i7_1_lut.init = 16'h5555;
    LUT4 inv_38_i6_1_lut (.A(xPre[5]), .Z(n280[5])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i6_1_lut.init = 16'h5555;
    LUT4 inv_38_i5_1_lut (.A(xPre[4]), .Z(n280[4])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i5_1_lut.init = 16'h5555;
    PFUMX i8311 (.BLUT(n11199), .ALUT(n11200), .C0(n12263), .Z(n11203));
    LUT4 i1327_4_lut (.A(n12228), .B(BUS_transferState[3]), .C(LOGIC_CLOCK_enable_26), 
         .D(n10846), .Z(LOGIC_CLOCK_enable_16)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(323[4] 373[11])
    defparam i1327_4_lut.init = 16'hcfc8;
    LUT4 i8597_3_lut_rep_193_4_lut (.A(\BUS_ADDR_INTERNAL[18]_derived_1 ), 
         .B(n1921), .C(n2129), .D(BUS_VALID_N_480), .Z(n12219)) /* synthesis lut_function=(A (B (C+!(D)))+!A (C+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[7:26])
    defparam i8597_3_lut_rep_193_4_lut.init = 16'hd0dd;
    LUT4 inv_38_i4_1_lut (.A(xPre[3]), .Z(n280[3])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i4_1_lut.init = 16'h5555;
    FD1P3DX xPre_681__i2 (.D(n37[2]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[2])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i2.GSR = "DISABLED";
    FD1P3DX xPre_681__i3 (.D(n37[3]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[3])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i3.GSR = "DISABLED";
    FD1P3DX xPre_681__i4 (.D(n37[4]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[4])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i4.GSR = "DISABLED";
    FD1P3DX xPre_681__i5 (.D(n37[5]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[5])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i5.GSR = "DISABLED";
    FD1P3DX xPre_681__i6 (.D(n37[6]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[6])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i6.GSR = "DISABLED";
    FD1P3DX xPre_681__i7 (.D(n37[7]), .SP(LOGIC_CLOCK_enable_167), .CK(LOGIC_CLOCK), 
            .CD(MATRIX_CURRROW_0_derived_5), .Q(xPre[7])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681__i7.GSR = "DISABLED";
    LUT4 inv_38_i3_1_lut (.A(xPre[2]), .Z(n280[2])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i3_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_159 (.A(n10309), .B(n11149), .C(Sprite_readData_15__N_417[12]), 
         .D(n12265), .Z(\MDM_data[12] )) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(49[8:16])
    defparam i1_4_lut_adj_159.init = 16'h5044;
    PFUMX i8312 (.BLUT(n11201), .ALUT(n11202), .C0(n12263), .Z(n11204));
    LUT4 inv_38_i2_1_lut (.A(xPre[1]), .Z(n280[1])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i2_1_lut.init = 16'h5555;
    PFUMX i8316 (.BLUT(n11206), .ALUT(n11207), .C0(n12263), .Z(Sprite_readData_15__N_417[5]));
    FD1P3DX currRowOffset_682__i1 (.D(n1[1]), .SP(LOGIC_CLOCK_enable_167), 
            .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), .Q(currRowOffset[1]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currRowOffset_682__i1.GSR = "DISABLED";
    PFUMX i8319 (.BLUT(n11209), .ALUT(n11210), .C0(n12263), .Z(Sprite_readData_15__N_417[6]));
    PFUMX i8322 (.BLUT(n11212), .ALUT(n11213), .C0(n12263), .Z(Sprite_readData_15__N_417[7]));
    LUT4 i1053_2_lut (.A(y[5]), .B(currRowOffset[0]), .Z(n162[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[48:59])
    defparam i1053_2_lut.init = 16'h6666;
    FD1P3AX currValue_i0_i1 (.D(BUS_data[1]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i1.GSR = "DISABLED";
    FD1P3AX currValue_i0_i2 (.D(BUS_data[2]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i2.GSR = "DISABLED";
    FD1P3AX currValue_i0_i3 (.D(BUS_data[3]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i3.GSR = "DISABLED";
    FD1P3AX currValue_i0_i4 (.D(BUS_data[4]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i4.GSR = "DISABLED";
    FD1P3AX currValue_i0_i5 (.D(BUS_data[5]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i5.GSR = "DISABLED";
    FD1P3AX currValue_i0_i6 (.D(BUS_data[6]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i6.GSR = "DISABLED";
    FD1P3AX currValue_i0_i7 (.D(BUS_data[7]), .SP(LOGIC_CLOCK_enable_175), 
            .CK(LOGIC_CLOCK), .Q(currValue[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=7, LSE_RCOL=35, LSE_LLINE=167, LSE_RLINE=167 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam currValue_i0_i7.GSR = "DISABLED";
    FD1P3DX currColor_683__i1 (.D(n12050), .SP(LOGIC_CLOCK_enable_178), 
            .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), .Q(currColor[1]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_683__i1.GSR = "DISABLED";
    FD1P3DX currColor_683__i2 (.D(n12049), .SP(LOGIC_CLOCK_enable_178), 
            .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), .Q(currColor[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_683__i2.GSR = "DISABLED";
    FD1P3DX currColor_683__i3 (.D(n12048), .SP(LOGIC_CLOCK_enable_178), 
            .CK(LOGIC_CLOCK), .CD(MATRIX_CURRROW_0_derived_5), .Q(currColor[3]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currColor_683__i3.GSR = "DISABLED";
    PFUMX i8327 (.BLUT(n11215), .ALUT(n11216), .C0(n12263), .Z(n11219));
    CCU2D xPre_681_add_4_9 (.A0(xPre[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10033), .S0(n37[7]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681_add_4_9.INIT0 = 16'hfaaa;
    defparam xPre_681_add_4_9.INIT1 = 16'h0000;
    defparam xPre_681_add_4_9.INJECT1_0 = "NO";
    defparam xPre_681_add_4_9.INJECT1_1 = "NO";
    LUT4 i7231_2_lut (.A(currRowOffset[1]), .B(currRowOffset[0]), .Z(n1[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i7231_2_lut.init = 16'h6666;
    CCU2D xPre_681_add_4_7 (.A0(xPre[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10032), .COUT(n10033), .S0(n37[5]), .S1(n37[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681_add_4_7.INIT0 = 16'hfaaa;
    defparam xPre_681_add_4_7.INIT1 = 16'hfaaa;
    defparam xPre_681_add_4_7.INJECT1_0 = "NO";
    defparam xPre_681_add_4_7.INJECT1_1 = "NO";
    PFUMX i8328 (.BLUT(n11217), .ALUT(n11218), .C0(n12263), .Z(n11220));
    LUT4 lastAddress_i1_i19_3_lut_3_lut_4_lut (.A(n12344), .B(n12304), .C(\lastAddress[18] ), 
         .D(SRAM_WE_N_704), .Z(n46)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C+!(D))) */ ;
    defparam lastAddress_i1_i19_3_lut_3_lut_4_lut.init = 16'hf0dd;
    LUT4 i7310_2_lut (.A(currAddress_17__N_488[8]), .B(y[1]), .Z(currAddress_17__N_488[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i7310_2_lut.init = 16'h6666;
    LUT4 i4753_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(n12304), .C(n2025), 
         .D(n12292), .Z(GR_WR_ADDR[1])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i4753_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_705_I_0_265_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12304), .C(n12292), .D(n13140), .Z(lastAddress_31__N_789)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_705_I_0_265_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 i4757_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(n12304), .C(n2025), 
         .D(n12272), .Z(GR_WR_ADDR[5])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i4757_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 i1_2_lut_2_lut_3_lut_3_lut_4_lut (.A(n12344), .B(n12304), .C(\BUS_addr[13] ), 
         .D(n13140), .Z(lastAddress_31__N_845)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam i1_2_lut_2_lut_3_lut_3_lut_4_lut.init = 16'h0f0d;
    LUT4 SRAM_WE_N_705_I_0_261_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12304), .C(n12272), .D(n13140), .Z(lastAddress_31__N_785)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_705_I_0_261_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 SRAM_WE_N_705_I_0_292_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12304), .C(n12288), .D(n13140), .Z(lastAddress_31__N_863)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam SRAM_WE_N_705_I_0_292_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 SRAM_WE_N_705_I_0_263_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12304), .C(n12287), .D(n13140), .Z(lastAddress_31__N_787)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_705_I_0_263_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5d5;
    LUT4 i4759_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(n12304), .C(n2025), 
         .D(n12288), .Z(GR_WR_ADDR[7])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i4759_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_705_I_0_259_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12304), .C(n12288), .D(n13140), .Z(lastAddress_31__N_783)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_705_I_0_259_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5d5;
    PFUMX i8332 (.BLUT(n11222), .ALUT(n11223), .C0(n12263), .Z(Sprite_readData_15__N_417[8]));
    LUT4 SRAM_WE_N_705_I_0_255_2_lut_2_lut_3_lut_3_lut_4_lut (.A(n12344), 
         .B(n12304), .C(\BUS_addr[11] ), .D(n13140), .Z(lastAddress_31__N_779)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam SRAM_WE_N_705_I_0_255_2_lut_2_lut_3_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 SRAM_WE_N_705_I_0_288_2_lut_2_lut_3_lut_3_lut_4_lut (.A(n12344), 
         .B(n12304), .C(\BUS_addr[11] ), .D(n13140), .Z(lastAddress_31__N_851)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam SRAM_WE_N_705_I_0_288_2_lut_2_lut_3_lut_3_lut_4_lut.init = 16'h0f0d;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), .B(n12304), 
         .C(n12272), .D(n13140), .Z(lastAddress_31__N_869)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0a08;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_160 (.A(n12344), .B(n12304), 
         .C(n12287), .D(n13140), .Z(lastAddress_31__N_875)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_160.init = 16'h0a08;
    LUT4 i4756_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(n12304), .C(n2025), 
         .D(n12278), .Z(GR_WR_ADDR[4])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i4756_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_161 (.A(n12344), .B(n12304), 
         .C(n12292), .D(n13140), .Z(lastAddress_31__N_881)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_161.init = 16'h0a08;
    LUT4 i4755_2_lut_3_lut_4_lut_4_lut (.A(n12344), .B(n12304), .C(n2025), 
         .D(n12287), .Z(GR_WR_ADDR[3])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C))) */ ;
    defparam i4755_2_lut_3_lut_4_lut_4_lut.init = 16'h0d05;
    LUT4 SRAM_WE_N_705_I_0_253_2_lut_2_lut_3_lut_3_lut_4_lut (.A(n12344), 
         .B(n12304), .C(\BUS_addr[13] ), .D(n13140), .Z(lastAddress_31__N_777)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam SRAM_WE_N_705_I_0_253_2_lut_2_lut_3_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i1_2_lut_2_lut_3_lut_3_lut_4_lut_adj_162 (.A(n12344), .B(n12304), 
         .C(\BUS_addr[14] ), .D(n13140), .Z(lastAddress_31__N_842)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam i1_2_lut_2_lut_3_lut_3_lut_4_lut_adj_162.init = 16'h0f0d;
    LUT4 SRAM_WE_N_705_I_0_252_2_lut_2_lut_3_lut_3_lut_4_lut (.A(n12344), 
         .B(n12304), .C(\BUS_addr[14] ), .D(n13140), .Z(lastAddress_31__N_776)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam SRAM_WE_N_705_I_0_252_2_lut_2_lut_3_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_163 (.A(n12344), .B(n12304), 
         .C(n12291), .D(n13140), .Z(lastAddress_31__N_857)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_163.init = 16'h0a08;
    LUT4 i4831_2_lut_rep_200_3_lut_3_lut_4_lut (.A(n12344), .B(n12304), 
         .C(n2025), .D(n13141), .Z(n12226)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (C (D)))) */ ;
    defparam i4831_2_lut_rep_200_3_lut_3_lut_4_lut.init = 16'h0dff;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_164 (.A(n12344), .B(n12304), 
         .C(n12278), .D(n13140), .Z(lastAddress_31__N_872)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut_adj_164.init = 16'h0a08;
    LUT4 SRAM_WE_N_705_I_0_262_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n12344), 
         .B(n12304), .C(n12278), .D(n13140), .Z(lastAddress_31__N_786)) /* synthesis lut_function=((B (C)+!B (C (D)))+!A) */ ;
    defparam SRAM_WE_N_705_I_0_262_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf5d5;
    PFUMX i8335 (.BLUT(n11225), .ALUT(n11226), .C0(n12263), .Z(Sprite_readData_15__N_417[9]));
    LUT4 i787_1_lut (.A(BUS_transferState[3]), .Z(GR_WR_CLK_N_689)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(315[3] 374[10])
    defparam i787_1_lut.init = 16'h5555;
    LUT4 i2_2_lut_rep_185_3_lut_4_lut (.A(n12331), .B(state[1]), .C(BUS_DONE), 
         .D(state[0]), .Z(LOGIC_CLOCK_enable_178)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_2_lut_rep_185_3_lut_4_lut.init = 16'h1000;
    PFUMX i8338 (.BLUT(n11228), .ALUT(n11229), .C0(n12263), .Z(Sprite_readData_15__N_417[12]));
    CCU2D xPre_681_add_4_5 (.A0(xPre[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10031), .COUT(n10032), .S0(n37[3]), .S1(n37[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681_add_4_5.INIT0 = 16'hfaaa;
    defparam xPre_681_add_4_5.INIT1 = 16'hfaaa;
    defparam xPre_681_add_4_5.INJECT1_0 = "NO";
    defparam xPre_681_add_4_5.INJECT1_1 = "NO";
    CCU2D xPre_681_add_4_3 (.A0(xPre[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(xPre[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10030), .COUT(n10031), .S0(n37[1]), .S1(n37[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681_add_4_3.INIT0 = 16'hfaaa;
    defparam xPre_681_add_4_3.INIT1 = 16'hfaaa;
    defparam xPre_681_add_4_3.INJECT1_0 = "NO";
    defparam xPre_681_add_4_3.INJECT1_1 = "NO";
    PFUMX i8341 (.BLUT(n11231), .ALUT(n11232), .C0(n12263), .Z(Sprite_readData_15__N_417[11]));
    PFUMX i8344 (.BLUT(n11234), .ALUT(n11235), .C0(n12263), .Z(Sprite_readData_15__N_417[13]));
    CCU2D xPre_681_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currRowOffset[0]), .B1(currRowOffset[1]), 
          .C1(xPre[0]), .D1(GND_net), .COUT(n10030), .S1(n37[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam xPre_681_add_4_1.INIT0 = 16'hF000;
    defparam xPre_681_add_4_1.INIT1 = 16'h7878;
    defparam xPre_681_add_4_1.INJECT1_0 = "NO";
    defparam xPre_681_add_4_1.INJECT1_1 = "NO";
    LUT4 i3_3_lut_4_lut_adj_165 (.A(n1184), .B(n12230), .C(BUS_DONE_OUT_N_627), 
         .D(n63), .Z(n8)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(323[4] 373[11])
    defparam i3_3_lut_4_lut_adj_165.init = 16'h0800;
    LUT4 BUS_DONE_OUT_I_45_2_lut_rep_202 (.A(BUS_DONE_OUT_N_626), .B(n2129), 
         .Z(n12228)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(355[11:65])
    defparam BUS_DONE_OUT_I_45_2_lut_rep_202.init = 16'h2222;
    LUT4 pwr_bdd_2_lut_rep_198_3_lut (.A(BUS_DONE_OUT_N_626), .B(n2129), 
         .C(n12157), .Z(n12224)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(355[11:65])
    defparam pwr_bdd_2_lut_rep_198_3_lut.init = 16'hfdfd;
    LUT4 i3_4_lut (.A(currColor[1]), .B(LOGIC_CLOCK_enable_178), .C(currColor[0]), 
         .D(n12343), .Z(LOGIC_CLOCK_enable_167)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i3_4_lut.init = 16'h0008;
    CCU2D add_431_19 (.A0(currAddress_17__N_488[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10029), .S0(currAddress[17]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_19.INIT0 = 16'h5aaa;
    defparam add_431_19.INIT1 = 16'h0000;
    defparam add_431_19.INJECT1_0 = "NO";
    defparam add_431_19.INJECT1_1 = "NO";
    PFUMX i8347 (.BLUT(n11237), .ALUT(n11238), .C0(n12263), .Z(Sprite_readData_15__N_417[10]));
    LUT4 i7_4_lut (.A(n13_adj_1297), .B(n11), .C(xPre[1]), .D(xPre[7]), 
         .Z(n15_adj_1298)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[8:20])
    defparam i7_4_lut.init = 16'hfeff;
    LUT4 i5_4_lut_adj_166 (.A(xPre[0]), .B(xPre[2]), .C(xPre[6]), .D(xPre[4]), 
         .Z(n13_adj_1297)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[8:20])
    defparam i5_4_lut_adj_166.init = 16'hfffe;
    LUT4 i3_2_lut (.A(xPre[3]), .B(xPre[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(250[8:20])
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i8730_2_lut (.A(n1627), .B(n1956), .Z(n11093)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(292[2] 295[36])
    defparam i8730_2_lut.init = 16'heeee;
    PFUMX i8220 (.BLUT(n11108), .ALUT(n11109), .C0(n12263), .Z(n11112));
    LUT4 i7229_1_lut (.A(currRowOffset[0]), .Z(n1[0])) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i7229_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(state[1]), .B(n8148), .C(state[0]), .Z(n10436)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i5630_3_lut (.A(state[4]), .B(n15_adj_1298), .C(state[2]), .Z(n8148)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i5630_3_lut.init = 16'h1a1a;
    PFUMX i8221 (.BLUT(n11110), .ALUT(n11111), .C0(n12263), .Z(n11113));
    CCU2D add_431_17 (.A0(currAddress_17__N_488[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_488[16]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n10028), .COUT(n10029), .S0(currAddress[15]), 
          .S1(currAddress[16]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_17.INIT0 = 16'h5aaa;
    defparam add_431_17.INIT1 = 16'h5aaa;
    defparam add_431_17.INJECT1_0 = "NO";
    defparam add_431_17.INJECT1_1 = "NO";
    CCU2D add_431_15 (.A0(currAddress_17__N_488[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_488[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n10027), .COUT(n10028), .S0(currAddress[13]), 
          .S1(currAddress[14]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_15.INIT0 = 16'h5aaa;
    defparam add_431_15.INIT1 = 16'h5aaa;
    defparam add_431_15.INJECT1_0 = "NO";
    defparam add_431_15.INJECT1_1 = "NO";
    PFUMX i8227 (.BLUT(n11115), .ALUT(n11116), .C0(n12263), .Z(n11119));
    LUT4 i8_4_lut (.A(n12276), .B(n11012), .C(n12274), .D(n12273), .Z(n18)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i8_4_lut.init = 16'h0010;
    LUT4 i8704_4_lut (.A(MATRIX_CURRROW[0]), .B(n12338), .C(state[4]), 
         .D(n11068), .Z(LOGIC_CLOCK_enable_1)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam i8704_4_lut.init = 16'h1000;
    LUT4 i8177_4_lut (.A(MATRIX_CURRROW[2]), .B(MATRIX_CURRROW[1]), .C(MATRIX_CURRROW[3]), 
         .D(MATRIX_CURRROW[4]), .Z(n11068)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8177_4_lut.init = 16'h8000;
    PFUMX i8228 (.BLUT(n11117), .ALUT(n11118), .C0(n12263), .Z(n11120));
    LUT4 i8153_2_lut (.A(\BUS_ADDR_INTERNAL[14] ), .B(\BUS_ADDR_INTERNAL[11] ), 
         .Z(n11052)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8153_2_lut.init = 16'heeee;
    PFUMX i8234 (.BLUT(n11122), .ALUT(n11123), .C0(n12263), .Z(n11126));
    LUT4 i4_4_lut_rep_208 (.A(n10350), .B(n8_adj_1299), .C(lastReadRow[0]), 
         .D(MATRIX_CURRROW[0]), .Z(MATRIX_CURRROW_0_derived_5)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[11:36])
    defparam i4_4_lut_rep_208.init = 16'hfeef;
    LUT4 i3_4_lut_adj_167 (.A(n12342), .B(n6), .C(lastReadRow[2]), .D(MATRIX_CURRROW[2]), 
         .Z(n8_adj_1299)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[11:36])
    defparam i3_4_lut_adj_167.init = 16'hedde;
    LUT4 lastReadRow_4__I_0_i10_1_lut_4_lut (.A(n10350), .B(n8_adj_1299), 
         .C(lastReadRow[0]), .D(MATRIX_CURRROW[0]), .Z(state_7__N_322)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[11:36])
    defparam lastReadRow_4__I_0_i10_1_lut_4_lut.init = 16'h0110;
    LUT4 i1_4_lut_adj_168 (.A(MATRIX_CURRROW[0]), .B(n10349), .C(lastReadRow[1]), 
         .D(MATRIX_CURRROW[1]), .Z(n6)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[11:36])
    defparam i1_4_lut_adj_168.init = 16'hedde;
    LUT4 i1_2_lut_3_lut_adj_169 (.A(n12232), .B(currRowOffset_lat[0]), .C(currRowOffset_lat[1]), 
         .Z(n3301)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_169.init = 16'h2020;
    LUT4 i1_4_lut_adj_170 (.A(n12327), .B(n19), .C(state[1]), .D(n160), 
         .Z(reset_N_670)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_170.init = 16'hcecc;
    LUT4 i1_4_lut_adj_171 (.A(reset), .B(state[1]), .C(n12331), .D(state[0]), 
         .Z(n19)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i1_4_lut_adj_171.init = 16'ha0a8;
    LUT4 i1_2_lut (.A(reset), .B(BUS_DONE), .Z(n160)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(34[8:13])
    defparam i1_2_lut.init = 16'heeee;
    PFUMX i8235 (.BLUT(n11124), .ALUT(n11125), .C0(n12263), .Z(n11127));
    LUT4 GR_WR_DOUT_9__I_0_i1_3_lut (.A(Sprite_readData[0]), .B(GR_WR_DOUT[0]), 
         .C(n1956), .Z(otherData[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(298[15:77])
    defparam GR_WR_DOUT_9__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 GR_WR_DOUT_9__I_0_i2_3_lut (.A(Sprite_readData[1]), .B(GR_WR_DOUT[1]), 
         .C(n1956), .Z(otherData[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(298[15:77])
    defparam GR_WR_DOUT_9__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 i1066_4_lut_3_lut_4_lut (.A(y[5]), .B(currRowOffset[0]), .C(y[6]), 
         .D(currRowOffset[1]), .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[48:59])
    defparam i1066_4_lut_3_lut_4_lut.init = 16'hf880;
    LUT4 i2_3_lut_4_lut (.A(y[5]), .B(currRowOffset[0]), .C(y[6]), .D(currRowOffset[1]), 
         .Z(n10348)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[48:59])
    defparam i2_3_lut_4_lut.init = 16'h8778;
    PFUMX i8241 (.BLUT(n11129), .ALUT(n11130), .C0(n12263), .Z(n11133));
    LUT4 i1_2_lut_3_lut_adj_172 (.A(y[5]), .B(currRowOffset[0]), .C(y[6]), 
         .Z(n4_adj_1294)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[48:59])
    defparam i1_2_lut_3_lut_adj_172.init = 16'h7878;
    LUT4 GR_WR_DOUT_9__I_0_i3_3_lut (.A(Sprite_readData[2]), .B(GR_WR_DOUT[2]), 
         .C(n1956), .Z(otherData[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(298[15:77])
    defparam GR_WR_DOUT_9__I_0_i3_3_lut.init = 16'hcaca;
    PFUMX i8242 (.BLUT(n11131), .ALUT(n11132), .C0(n12263), .Z(n11134));
    LUT4 i8697_2_lut_4_lut_4_lut (.A(n12244), .B(n12218), .C(n12269), 
         .D(n12265), .Z(n3242)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i8697_2_lut_4_lut_4_lut.init = 16'h0010;
    CCU2D add_431_13 (.A0(currAddress_17__N_488[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_488[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n10026), .COUT(n10027), .S0(currAddress[11]), 
          .S1(currAddress[12]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_13.INIT0 = 16'h5aaa;
    defparam add_431_13.INIT1 = 16'h5aaa;
    defparam add_431_13.INJECT1_0 = "NO";
    defparam add_431_13.INJECT1_1 = "NO";
    CCU2D add_431_11 (.A0(currAddress_17__N_488[9]), .B0(currAddress_17__N_506[9]), 
          .C0(GND_net), .D0(GND_net), .A1(currAddress_17__N_488[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10025), .COUT(n10026), 
          .S0(currAddress[9]), .S1(currAddress[10]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_11.INIT0 = 16'h5666;
    defparam add_431_11.INIT1 = 16'h5aaa;
    defparam add_431_11.INJECT1_0 = "NO";
    defparam add_431_11.INJECT1_1 = "NO";
    LUT4 i2210_4_lut (.A(n12344), .B(n12304), .C(n13158), .D(n12280), 
         .Z(BUS_VALID_N_480)) /* synthesis lut_function=((B ((D)+!C))+!A) */ ;
    defparam i2210_4_lut.init = 16'hdd5d;
    LUT4 GR_WR_DOUT_9__I_0_i4_3_lut (.A(Sprite_readData[3]), .B(GR_WR_DOUT[3]), 
         .C(n1956), .Z(otherData[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(298[15:77])
    defparam GR_WR_DOUT_9__I_0_i4_3_lut.init = 16'hcaca;
    PFUMX i8436 (.BLUT(n11324), .ALUT(n11325), .C0(n12263), .Z(n11328));
    LUT4 i8710_2_lut_4_lut_4_lut (.A(n12244), .B(n12218), .C(n12269), 
         .D(n12292), .Z(n3137)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i8710_2_lut_4_lut_4_lut.init = 16'h0001;
    CCU2D add_431_9 (.A0(currAddress_17__N_506[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_488[8]), .B1(currAddress_17__N_506[8]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10024), .COUT(n10025), .S0(currAddress[7]), 
          .S1(currAddress[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_9.INIT0 = 16'hfaaa;
    defparam add_431_9.INIT1 = 16'h5666;
    defparam add_431_9.INJECT1_0 = "NO";
    defparam add_431_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_173 (.A(state[0]), .B(BUS_DONE), .C(MATRIX_CURRROW_0_derived_5), 
         .D(n12297), .Z(LOGIC_CLOCK_enable_175)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_173.init = 16'h0008;
    LUT4 mux_553_i1_3_lut_4_lut (.A(n12292), .B(n12344), .C(latchMode[0]), 
         .D(n2266), .Z(n2372[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam mux_553_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_6_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[6]), .D(n11205), .Z(Sprite_readData[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_6_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_7_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[7]), .D(n11330), .Z(Sprite_readData[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_7_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_9_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[9]), .D(n11128), .Z(Sprite_readData[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_9_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i25_3_lut_4_lut (.A(n12292), .B(n12344), .C(Sprite_readData_15__N_417[15]), 
         .D(n11170), .Z(n12_adj_1295)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam i25_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_8_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[8]), .D(n11121), .Z(Sprite_readData[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_8_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_0_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[0]), .D(n11192), .Z(Sprite_readData[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_0_i3_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i8437 (.BLUT(n11326), .ALUT(n11327), .C0(n12263), .Z(n11329));
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_4_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[4]), .D(n11337), .Z(Sprite_readData[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_4_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_5_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[5]), .D(n11221), .Z(Sprite_readData[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_5_i3_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i8248 (.BLUT(n11136), .ALUT(n11137), .C0(n12263), .Z(n11140));
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_3_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[3]), .D(n11100), .Z(Sprite_readData[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_3_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i2_3_lut_rep_204_4_lut (.A(n12292), .B(n12344), .C(n10855), .D(n12277), 
         .Z(n12230)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam i2_3_lut_rep_204_4_lut.init = 16'hfbff;
    LUT4 lastAddress_i1_i2_3_lut_3_lut_4_lut (.A(n12292), .B(n12344), .C(\lastAddress[1] ), 
         .D(SRAM_WE_N_704), .Z(n63_adj_34)) /* synthesis lut_function=(A (C+!(D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam lastAddress_i1_i2_3_lut_3_lut_4_lut.init = 16'hf0bb;
    LUT4 mux_553_i2_3_lut_4_lut (.A(n12292), .B(n12344), .C(latchMode[1]), 
         .D(n2265), .Z(n2372[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam mux_553_i2_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i8443 (.BLUT(n11331), .ALUT(n11332), .C0(n12263), .Z(n11335));
    LUT4 mux_553_i3_3_lut_4_lut (.A(n12292), .B(n12344), .C(latchMode[2]), 
         .D(n2264), .Z(n2372[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam mux_553_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_553_i4_3_lut_4_lut (.A(n12292), .B(n12344), .C(latchMode[3]), 
         .D(n2263), .Z(n2372[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam mux_553_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_2_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[2]), .D(n11107), .Z(Sprite_readData[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_2_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 BUS_ADDR_IN_1__I_0_413_Mux_1_i3_3_lut_4_lut (.A(n12292), .B(n12344), 
         .C(Sprite_readData_15__N_417[1]), .D(n11114), .Z(Sprite_readData[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(167[7:35])
    defparam BUS_ADDR_IN_1__I_0_413_Mux_1_i3_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i8444 (.BLUT(n11333), .ALUT(n11334), .C0(n12263), .Z(n11336));
    LUT4 i2_3_lut_rep_206_4_lut (.A(n12331), .B(state[0]), .C(MATRIX_CURRROW_0_derived_5), 
         .D(state[1]), .Z(n12232)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_rep_206_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_174 (.A(n12331), .B(state[0]), .C(n11_adj_1301), 
         .D(state[1]), .Z(n10870)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_174.init = 16'h0400;
    PFUMX i8249 (.BLUT(n11138), .ALUT(n11139), .C0(n12263), .Z(n11141));
    LUT4 i1_2_lut_rep_305 (.A(state[2]), .B(state[4]), .Z(n12331)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i1_2_lut_rep_305.init = 16'heeee;
    LUT4 i54_2_lut_3_lut (.A(state[2]), .B(state[4]), .C(BUS_DONE), .Z(n54)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i54_2_lut_3_lut.init = 16'h0101;
    PFUMX i8255 (.BLUT(n11143), .ALUT(n11144), .C0(n12263), .Z(n11147));
    LUT4 i8107_2_lut_rep_271_3_lut (.A(state[2]), .B(state[4]), .C(state[1]), 
         .Z(n12297)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i8107_2_lut_rep_271_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut_rep_268_3_lut_4_lut (.A(state[2]), .B(state[4]), .C(state[1]), 
         .D(state[0]), .Z(LOGIC_CLOCK_N_116_enable_20)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i2_2_lut_rep_268_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_301_3_lut (.A(state[2]), .B(state[4]), .C(state[0]), 
         .Z(n12327)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(53[9:14])
    defparam i1_2_lut_rep_301_3_lut.init = 16'h1010;
    CCU2D add_431_7 (.A0(currAddress_17__N_506[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_506[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10023), .COUT(n10024), .S0(currAddress[5]), 
          .S1(currAddress[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_7.INIT0 = 16'hfaaa;
    defparam add_431_7.INIT1 = 16'hfaaa;
    defparam add_431_7.INJECT1_0 = "NO";
    defparam add_431_7.INJECT1_1 = "NO";
    PFUMX i8256 (.BLUT(n11145), .ALUT(n11146), .C0(n12263), .Z(n11148));
    LUT4 offsetLatchClock_I_0_4_lut (.A(LOGIC_CLOCK), .B(latchForce), .C(n10893), 
         .D(n9), .Z(offsetLatchClockOrd)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(169[25:55])
    defparam offsetLatchClock_I_0_4_lut.init = 16'hfcee;
    LUT4 i1_3_lut (.A(latchMode[1]), .B(frameEndClock), .C(latchMode[0]), 
         .Z(n10893)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut.init = 16'h0808;
    LUT4 i2_4_lut_adj_175 (.A(latchMode[1]), .B(latchMode[2]), .C(latchMode[0]), 
         .D(latchMode[3]), .Z(n9)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+((D)+!C)))) */ ;
    defparam i2_4_lut_adj_175.init = 16'h0012;
    CCU2D add_431_5 (.A0(currColor[3]), .B0(currAddress_17__N_506[3]), .C0(GND_net), 
          .D0(GND_net), .A1(currAddress_17__N_506[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10022), .COUT(n10023), .S0(currAddress[3]), 
          .S1(currAddress[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_5.INIT0 = 16'h5666;
    defparam add_431_5.INIT1 = 16'hfaaa;
    defparam add_431_5.INJECT1_0 = "NO";
    defparam add_431_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_176 (.A(state[2]), .B(state[1]), .C(n21), .D(n24), 
         .Z(n10478)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_176.init = 16'h7350;
    CCU2D add_431_3 (.A0(currColor[1]), .B0(currAddress_17__N_506[1]), .C0(GND_net), 
          .D0(GND_net), .A1(currColor[2]), .B1(currAddress_17__N_506[2]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10021), .COUT(n10022), .S0(currAddress[1]), 
          .S1(currAddress[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_3.INIT0 = 16'h5666;
    defparam add_431_3.INIT1 = 16'h5666;
    defparam add_431_3.INJECT1_0 = "NO";
    defparam add_431_3.INJECT1_1 = "NO";
    CCU2D add_7182_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10204), 
          .S0(n2025));
    defparam add_7182_cout.INIT0 = 16'h0000;
    defparam add_7182_cout.INIT1 = 16'h0000;
    defparam add_7182_cout.INJECT1_0 = "NO";
    defparam add_7182_cout.INJECT1_1 = "NO";
    CCU2D add_7182_11 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n10203), .COUT(n10204));
    defparam add_7182_11.INIT0 = 16'heeee;
    defparam add_7182_11.INIT1 = 16'heeee;
    defparam add_7182_11.INJECT1_0 = "NO";
    defparam add_7182_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_177 (.A(state[4]), .B(n11060), .C(state[1]), .D(n11_adj_1301), 
         .Z(n21)) /* synthesis lut_function=(!(A (B)+!A !((C (D))+!B))) */ ;
    defparam i1_4_lut_adj_177.init = 16'h7333;
    LUT4 i8170_4_lut (.A(state[0]), .B(state[1]), .C(state[4]), .D(n12332), 
         .Z(n11060)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i8170_4_lut.init = 16'hfbfa;
    CCU2D add_431_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(xPre[0]), .B1(xOffset[0]), .C1(currColor[0]), .D1(GND_net), 
          .COUT(n10021), .S1(currAddress[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(166[47:168])
    defparam add_431_1.INIT0 = 16'hF000;
    defparam add_431_1.INIT1 = 16'h9696;
    defparam add_431_1.INJECT1_0 = "NO";
    defparam add_431_1.INJECT1_1 = "NO";
    CCU2D add_7182_9 (.A0(n13158), .B0(n12344), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), 
          .D1(n12309), .CIN(n10202), .COUT(n10203));
    defparam add_7182_9.INIT0 = 16'h8888;
    defparam add_7182_9.INIT1 = 16'hff20;
    defparam add_7182_9.INJECT1_0 = "NO";
    defparam add_7182_9.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_178 (.A(currColor_lat[0]), .B(currRowOffset_lat[1]), 
         .C(currRowOffset_lat[0]), .D(n10888), .Z(n11_adj_1301)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i3_4_lut_adj_178.init = 16'hffbf;
    LUT4 i2_3_lut_rep_312 (.A(state[2]), .B(state[0]), .C(state[1]), .Z(n12338)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam i2_3_lut_rep_312.init = 16'hfefe;
    LUT4 i2_3_lut_adj_179 (.A(currColor_lat[3]), .B(currColor_lat[1]), .C(currColor_lat[2]), 
         .Z(n10888)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i2_3_lut_adj_179.init = 16'hfbfb;
    LUT4 i8584_2_lut_2_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(MATRIX_CURRROW_0_derived_5), .Z(LOGIC_CLOCK_enable_6)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam i8584_2_lut_2_lut_4_lut.init = 16'h0001;
    LUT4 inv_38_i1_1_lut (.A(xPre[0]), .Z(n280[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(207[36:55])
    defparam inv_38_i1_1_lut.init = 16'h5555;
    LUT4 i8632_2_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(state[4]), .Z(n10852)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(183[3] 268[10])
    defparam i8632_2_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_180 (.A(n12220), .B(WRITE_DONE), .C(n10), .D(WRITE_DONE_adj_35), 
         .Z(BUS_DONE)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_180.init = 16'hfffe;
    LUT4 i1_3_lut_3_lut (.A(state[4]), .B(n15_adj_1298), .C(state[2]), 
         .Z(n14)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h4040;
    LUT4 i8123_2_lut_rep_317 (.A(currColor[3]), .B(currColor[2]), .Z(n12343)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8123_2_lut_rep_317.init = 16'heeee;
    LUT4 i4_4_lut (.A(n7), .B(BUS_DONE_OVERRIDE), .C(\BUS_ADDR_INTERNAL[18]_derived_1 ), 
         .D(BUS_DONE_INTERNAL), .Z(n10)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i4_4_lut.init = 16'hefee;
    LUT4 currColor_1__bdd_4_lut (.A(currColor[1]), .B(currColor[3]), .C(currColor[2]), 
         .D(currColor[0]), .Z(n12048)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B))) */ ;
    defparam currColor_1__bdd_4_lut.init = 16'h6ccc;
    LUT4 n11010_bdd_3_lut_4_lut (.A(currColor[3]), .B(currColor[2]), .C(currColor[0]), 
         .D(currColor[1]), .Z(n12050)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam n11010_bdd_3_lut_4_lut.init = 16'h0ef0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_181 (.A(currColor[3]), .B(currColor[2]), 
         .C(currColor[0]), .D(currColor[1]), .Z(n27[0])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_181.init = 16'h0e0f;
    CCU2D add_7182_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n13150), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16]_adj_19 ), 
          .D1(n13151), .CIN(n10201), .COUT(n10202));
    defparam add_7182_7.INIT0 = 16'h00ae;
    defparam add_7182_7.INIT1 = 16'h00ae;
    defparam add_7182_7.INJECT1_0 = "NO";
    defparam add_7182_7.INJECT1_1 = "NO";
    GammaRam GRam (.\BUS_data[9] (BUS_data[9]), .GND_net(GND_net), .GR_WR_ADDR({GR_WR_ADDR[7], 
            \GR_WR_ADDR[6] , GR_WR_ADDR[5:3], \GR_WR_ADDR[2] , GR_WR_ADDR[1], 
            \GR_WR_ADDR[0] }), .currValue({currValue}), .GR_WR_CLK(GR_WR_CLK), 
            .LOGIC_CLOCK_N_116(LOGIC_CLOCK_N_116), .VCC_net(VCC_net), .n13141(n13141), 
            .GR_WR_DOUT({GR_WR_DOUT[9:8], \GR_WR_DOUT[7] , \GR_WR_DOUT[6] , 
            \GR_WR_DOUT[5] , \GR_WR_DOUT[4] , GR_WR_DOUT[3:0]}), .GR_RE_DOUT({GR_RE_DOUT}), 
            .\BUS_data[8] (BUS_data[8]), .\BUS_data[7] (BUS_data[7]), .\BUS_data[6] (BUS_data[6]), 
            .\BUS_data[5] (BUS_data[5]), .\BUS_data[4] (BUS_data[4]), .\BUS_data[3] (BUS_data[3]), 
            .\BUS_data[2] (BUS_data[2]), .\BUS_data[1] (BUS_data[1]), .\BUS_data[0] (BUS_data[0])) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(381[8:16])
    
endmodule
//
// Verilog Description of module GammaRam
//

module GammaRam (\BUS_data[9] , GND_net, GR_WR_ADDR, currValue, GR_WR_CLK, 
            LOGIC_CLOCK_N_116, VCC_net, n13141, GR_WR_DOUT, GR_RE_DOUT, 
            \BUS_data[8] , \BUS_data[7] , \BUS_data[6] , \BUS_data[5] , 
            \BUS_data[4] , \BUS_data[3] , \BUS_data[2] , \BUS_data[1] , 
            \BUS_data[0] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input \BUS_data[9] ;
    input GND_net;
    input [7:0]GR_WR_ADDR;
    input [7:0]currValue;
    input GR_WR_CLK;
    input LOGIC_CLOCK_N_116;
    input VCC_net;
    input n13141;
    output [9:0]GR_WR_DOUT;
    output [9:0]GR_RE_DOUT;
    input \BUS_data[8] ;
    input \BUS_data[7] ;
    input \BUS_data[6] ;
    input \BUS_data[5] ;
    input \BUS_data[4] ;
    input \BUS_data[3] ;
    input \BUS_data[2] ;
    input \BUS_data[1] ;
    input \BUS_data[0] ;
    
    wire GR_WR_CLK /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(138[9:18])
    wire LOGIC_CLOCK_N_116 /* synthesis is_clock=1, is_inv_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(73[9:17])
    
    DP8KC GammaRam_0_1_0 (.DIA0(\BUS_data[9] ), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(VCC_net), .ADA1(GND_net), 
          .ADA2(GND_net), .ADA3(GR_WR_ADDR[0]), .ADA4(GR_WR_ADDR[1]), 
          .ADA5(GR_WR_ADDR[2]), .ADA6(GR_WR_ADDR[3]), .ADA7(GR_WR_ADDR[4]), 
          .ADA8(GR_WR_ADDR[5]), .ADA9(GR_WR_ADDR[6]), .ADA10(GR_WR_ADDR[7]), 
          .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), 
          .CLKA(GR_WR_CLK), .WEA(n13141), .CSA0(GND_net), .CSA1(GND_net), 
          .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
          .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
          .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), 
          .ADB1(GND_net), .ADB2(GND_net), .ADB3(currValue[0]), .ADB4(currValue[1]), 
          .ADB5(currValue[2]), .ADB6(currValue[3]), .ADB7(currValue[4]), 
          .ADB8(currValue[5]), .ADB9(currValue[6]), .ADB10(currValue[7]), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), 
          .CLKB(LOGIC_CLOCK_N_116), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(GND_net), .DOA0(GR_WR_DOUT[9]), .DOB0(GR_RE_DOUT[9])) /* synthesis MEM_LPC_FILE="GammaRam.lpc", MEM_INIT_FILE="gammadefault.mem", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=16, LSE_LLINE=381, LSE_RLINE=381 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(381[8:16])
    defparam GammaRam_0_1_0.DATA_WIDTH_A = 9;
    defparam GammaRam_0_1_0.DATA_WIDTH_B = 9;
    defparam GammaRam_0_1_0.REGMODE_A = "NOREG";
    defparam GammaRam_0_1_0.REGMODE_B = "NOREG";
    defparam GammaRam_0_1_0.CSDECODE_A = "0b000";
    defparam GammaRam_0_1_0.CSDECODE_B = "0b000";
    defparam GammaRam_0_1_0.WRITEMODE_A = "NORMAL";
    defparam GammaRam_0_1_0.WRITEMODE_B = "NORMAL";
    defparam GammaRam_0_1_0.GSR = "ENABLED";
    defparam GammaRam_0_1_0.RESETMODE = "ASYNC";
    defparam GammaRam_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam GammaRam_0_1_0.INIT_DATA = "STATIC";
    defparam GammaRam_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_04 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_05 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_06 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_07 = "0x00201002010020100201002010020100201002010020100201002010020100201002010020100201";
    defparam GammaRam_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC GammaRam_0_0_1 (.DIA0(\BUS_data[0] ), .DIA1(\BUS_data[1] ), .DIA2(\BUS_data[2] ), 
          .DIA3(\BUS_data[3] ), .DIA4(\BUS_data[4] ), .DIA5(\BUS_data[5] ), 
          .DIA6(\BUS_data[6] ), .DIA7(\BUS_data[7] ), .DIA8(\BUS_data[8] ), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(GR_WR_ADDR[0]), 
          .ADA4(GR_WR_ADDR[1]), .ADA5(GR_WR_ADDR[2]), .ADA6(GR_WR_ADDR[3]), 
          .ADA7(GR_WR_ADDR[4]), .ADA8(GR_WR_ADDR[5]), .ADA9(GR_WR_ADDR[6]), 
          .ADA10(GR_WR_ADDR[7]), .ADA11(GND_net), .ADA12(GND_net), .CEA(VCC_net), 
          .OCEA(VCC_net), .CLKA(GR_WR_CLK), .WEA(n13141), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(VCC_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(currValue[0]), 
          .ADB4(currValue[1]), .ADB5(currValue[2]), .ADB6(currValue[3]), 
          .ADB7(currValue[4]), .ADB8(currValue[5]), .ADB9(currValue[6]), 
          .ADB10(currValue[7]), .ADB11(GND_net), .ADB12(GND_net), .CEB(VCC_net), 
          .OCEB(VCC_net), .CLKB(LOGIC_CLOCK_N_116), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOA0(GR_WR_DOUT[0]), 
          .DOA1(GR_WR_DOUT[1]), .DOA2(GR_WR_DOUT[2]), .DOA3(GR_WR_DOUT[3]), 
          .DOA4(GR_WR_DOUT[4]), .DOA5(GR_WR_DOUT[5]), .DOA6(GR_WR_DOUT[6]), 
          .DOA7(GR_WR_DOUT[7]), .DOA8(GR_WR_DOUT[8]), .DOB0(GR_RE_DOUT[0]), 
          .DOB1(GR_RE_DOUT[1]), .DOB2(GR_RE_DOUT[2]), .DOB3(GR_RE_DOUT[3]), 
          .DOB4(GR_RE_DOUT[4]), .DOB5(GR_RE_DOUT[5]), .DOB6(GR_RE_DOUT[6]), 
          .DOB7(GR_RE_DOUT[7]), .DOB8(GR_RE_DOUT[8])) /* synthesis MEM_LPC_FILE="GammaRam.lpc", MEM_INIT_FILE="gammadefault.mem", syn_instantiated=1, LSE_LINE_FILE_ID=26, LSE_LCOL=8, LSE_RCOL=16, LSE_LLINE=381, LSE_RLINE=381 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixbushandler.vhd(381[8:16])
    defparam GammaRam_0_0_1.DATA_WIDTH_A = 9;
    defparam GammaRam_0_0_1.DATA_WIDTH_B = 9;
    defparam GammaRam_0_0_1.REGMODE_A = "NOREG";
    defparam GammaRam_0_0_1.REGMODE_B = "NOREG";
    defparam GammaRam_0_0_1.CSDECODE_A = "0b000";
    defparam GammaRam_0_0_1.CSDECODE_B = "0b000";
    defparam GammaRam_0_0_1.WRITEMODE_A = "NORMAL";
    defparam GammaRam_0_0_1.WRITEMODE_B = "NORMAL";
    defparam GammaRam_0_0_1.GSR = "ENABLED";
    defparam GammaRam_0_0_1.RESETMODE = "ASYNC";
    defparam GammaRam_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam GammaRam_0_0_1.INIT_DATA = "STATIC";
    defparam GammaRam_0_0_1.INITVAL_00 = "0x0F8780E8700D8680C8600B8580A85009848088400783806830058280482003818028100180800800";
    defparam GammaRam_0_0_1.INITVAL_01 = "0x1F8F81E8F01D8E81C8E01B8D81A8D0198C8188C0178B8168B0158A8148A013898128901188810880";
    defparam GammaRam_0_0_1.INITVAL_02 = "0x2F9782E9702D9682C9602B9582A95029948289402793826930259282492023918229102190820900";
    defparam GammaRam_0_0_1.INITVAL_03 = "0x3F9F83E9F03D9E83C9E03B9D83A9D0399C8389C0379B8369B0359A8349A033998329903198830980";
    defparam GammaRam_0_0_1.INITVAL_04 = "0x0F8780E8700D8680C8600B8580A85009848088400783806830058280482003818028100180800800";
    defparam GammaRam_0_0_1.INITVAL_05 = "0x1F8F81E8F01D8E81C8E01B8D81A8D0198C8188C0178B8168B0158A8148A013898128901188810880";
    defparam GammaRam_0_0_1.INITVAL_06 = "0x2F9782E9702D9682C9602B9582A95029948289402793826930259282492023918229102190820900";
    defparam GammaRam_0_0_1.INITVAL_07 = "0x3F9F83E9F03D9E83C9E03B9D83A9D0399C8389C0379B8369B0359A8349A033998329903198830980";
    defparam GammaRam_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam GammaRam_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module PIC
//

module PIC (GND_net, PIC_ADDR_IN_c_15, PIC_ADDR_IN_c_14, PIC_ADDR_IN_c_13, 
            PIC_ADDR_IN_c_12, state, LOGIC_CLOCK, \BUS_data[0] , \BUS_ADDR_INTERNAL[0] , 
            PIC_ADDR_IN_c_0, \BUS_req[2] , WRITE_DONE, transferMode_3__N_1115, 
            n13160, PIC_ADDR_IN_c_1, PIC_ADDR_IN_c_2, PIC_ADDR_IN_c_3, 
            PIC_ADDR_IN_c_4, PIC_ADDR_IN_c_5, PIC_ADDR_IN_c_6, PIC_ADDR_IN_c_7, 
            PIC_ADDR_IN_c_8, PIC_ADDR_IN_c_9, PIC_ADDR_IN_c_10, PIC_ADDR_IN_c_11, 
            PIC_ADDR_IN_c_16, PIC_ADDR_IN_c_17, PIC_ADDR_IN_c_18, n11758, 
            n5045, n12252, n12263, n87, BUS_VALID_N_1118, \BUS_currGrantID[0] , 
            \BUS_currGrantID[1] , n13158, n12344, \BUS_ADDR_INTERNAL[18] , 
            n12309, \BUS_ADDR_INTERNAL[15] , n13150, \BUS_ADDR_INTERNAL[16] , 
            n13151, \BUS_ADDR_INTERNAL[13] , n13155, \BUS_ADDR_INTERNAL[14] , 
            n13157, \BUS_ADDR_INTERNAL[11] , n13156, \BUS_ADDR_INTERNAL[12] , 
            n13142, \BUS_ADDR_INTERNAL[9] , n13144, \BUS_ADDR_INTERNAL[10] , 
            n13143, \BUS_ADDR_INTERNAL[8] , n13154, PIC_DATA_IN_out_15, 
            PIC_DATA_IN_out_13, PIC_DATA_IN_out_14, PIC_DATA_IN_out_11, 
            PIC_DATA_IN_out_12, PIC_DATA_IN_out_9, PIC_DATA_IN_out_10, 
            PIC_DATA_IN_out_8, PIC_READY_c, BUS_DIRECTION_INTERNAL, n2198, 
            \BUS_data[1] , \BUS_data[2] , \BUS_data[3] , \BUS_ADDR_INTERNAL[1] , 
            \BUS_ADDR_INTERNAL[2] , \BUS_ADDR_INTERNAL[3] , \BUS_ADDR_INTERNAL[4] , 
            \BUS_ADDR_INTERNAL[5] , \BUS_ADDR_INTERNAL[6] , \BUS_ADDR_INTERNAL[7] , 
            \BUS_ADDR_INTERNAL[8]_adj_1 , \BUS_ADDR_INTERNAL[9]_adj_2 , 
            \BUS_ADDR_INTERNAL[10]_adj_3 , \BUS_ADDR_INTERNAL[11]_adj_4 , 
            \BUS_ADDR_INTERNAL[12]_adj_5 , \BUS_ADDR_INTERNAL[13]_adj_6 , 
            \BUS_ADDR_INTERNAL[14]_adj_7 , \BUS_ADDR_INTERNAL[15]_adj_8 , 
            \BUS_ADDR_INTERNAL[16]_adj_9 , \BUS_ADDR_INTERNAL[17] , PIC_DATA_IN_out_3, 
            PIC_WE_IN_c, PIC_DATA_IN_out_6, n12276, n12274, n12291, 
            \BUS_ADDR_INTERNAL[5]_adj_10 , n12272, \BUS_ADDR_INTERNAL[6]_adj_11 , 
            n12289, \BUS_ADDR_INTERNAL[7]_adj_12 , n12288, PIC_DATA_IN_out_5, 
            PIC_DATA_IN_out_7, \BUS_ADDR_INTERNAL[3]_adj_13 , n12287, 
            n12290, \BUS_data[4] , \BUS_data[5] , \BUS_data[6] , \BUS_data[7] , 
            \BUS_ADDR_INTERNAL[1]_adj_14 , n12292, \writeData[4] , \writeData[5] , 
            \writeData[6] , \writeData[7] , n12280, n1921, n12222, 
            n2025, LOGIC_CLOCK_enable_26, \BUS_ADDR_INTERNAL[2]_adj_15 , 
            n12279, \BUS_ADDR_INTERNAL[4]_adj_16 , n12278, n13147, \state[7] , 
            \state_7__N_1050[7] , n12273, n13145, n13146, n13148, 
            n13153, n13149, n13152, \BUS_ADDR_INTERNAL[0]_adj_17 , n12299, 
            PIC_DATA_IN_out_1, PIC_DATA_IN_out_2, PIC_DATA_IN_out_4, n12223, 
            n13141, n11485, n12219, LOGIC_CLOCK_enable_48, n7167, 
            n12213, n12314, \BUS_DATA_INTERNAL[2] , n6, \BUS_currGrantID_3__N_72[0] , 
            \BUS_currGrantID_3__N_72[1] , n12352, n71, PIC_OE_c, n12312, 
            n12214, n12324, PIC_DATA_IN_out_0, n12212, n12348, n13139, 
            n6_adj_18, \BUS_DATA_INTERNAL[1] , n10895, n69, n1184, 
            BUS_currGrantID_3__N_54, BUS_DONE, \BUS_DATA_INTERNAL[0] , 
            n12250, n12217, \PIC_data[9] , \PIC_data[11] , \PIC_data[10] , 
            n100, \PIC_data[12] , \PIC_data[8] , \PIC_data[13] , \PIC_data[14] , 
            SRAM_WE_N_704, \lastAddress[4] , n60, n10904, \lastAddress[7] , 
            n57, \lastAddress[3] , n61, \lastAddress[17] , n47, n13140, 
            n12304, lastAddress_31__N_833, lastAddress_31__N_773, n9924, 
            BUS_DONE_OUT_N_626, \BUS_DATA_INTERNAL[3] , n12332, n10976, 
            n11012);
    input GND_net;
    input PIC_ADDR_IN_c_15;
    input PIC_ADDR_IN_c_14;
    input PIC_ADDR_IN_c_13;
    input PIC_ADDR_IN_c_12;
    output [7:0]state;
    input LOGIC_CLOCK;
    input \BUS_data[0] ;
    output \BUS_ADDR_INTERNAL[0] ;
    input PIC_ADDR_IN_c_0;
    output \BUS_req[2] ;
    output WRITE_DONE;
    input transferMode_3__N_1115;
    input n13160;
    input PIC_ADDR_IN_c_1;
    input PIC_ADDR_IN_c_2;
    input PIC_ADDR_IN_c_3;
    input PIC_ADDR_IN_c_4;
    input PIC_ADDR_IN_c_5;
    input PIC_ADDR_IN_c_6;
    input PIC_ADDR_IN_c_7;
    input PIC_ADDR_IN_c_8;
    input PIC_ADDR_IN_c_9;
    input PIC_ADDR_IN_c_10;
    input PIC_ADDR_IN_c_11;
    input PIC_ADDR_IN_c_16;
    input PIC_ADDR_IN_c_17;
    input PIC_ADDR_IN_c_18;
    input n11758;
    input n5045;
    input n12252;
    input n12263;
    output n87;
    output BUS_VALID_N_1118;
    input \BUS_currGrantID[0] ;
    input \BUS_currGrantID[1] ;
    input n13158;
    input n12344;
    output \BUS_ADDR_INTERNAL[18] ;
    input n12309;
    input \BUS_ADDR_INTERNAL[15] ;
    input n13150;
    input \BUS_ADDR_INTERNAL[16] ;
    input n13151;
    input \BUS_ADDR_INTERNAL[13] ;
    input n13155;
    input \BUS_ADDR_INTERNAL[14] ;
    input n13157;
    input \BUS_ADDR_INTERNAL[11] ;
    input n13156;
    input \BUS_ADDR_INTERNAL[12] ;
    input n13142;
    input \BUS_ADDR_INTERNAL[9] ;
    input n13144;
    input \BUS_ADDR_INTERNAL[10] ;
    input n13143;
    input \BUS_ADDR_INTERNAL[8] ;
    input n13154;
    input PIC_DATA_IN_out_15;
    input PIC_DATA_IN_out_13;
    input PIC_DATA_IN_out_14;
    input PIC_DATA_IN_out_11;
    input PIC_DATA_IN_out_12;
    input PIC_DATA_IN_out_9;
    input PIC_DATA_IN_out_10;
    input PIC_DATA_IN_out_8;
    output PIC_READY_c;
    output BUS_DIRECTION_INTERNAL;
    output n2198;
    input \BUS_data[1] ;
    input \BUS_data[2] ;
    input \BUS_data[3] ;
    output \BUS_ADDR_INTERNAL[1] ;
    output \BUS_ADDR_INTERNAL[2] ;
    output \BUS_ADDR_INTERNAL[3] ;
    output \BUS_ADDR_INTERNAL[4] ;
    output \BUS_ADDR_INTERNAL[5] ;
    output \BUS_ADDR_INTERNAL[6] ;
    output \BUS_ADDR_INTERNAL[7] ;
    output \BUS_ADDR_INTERNAL[8]_adj_1 ;
    output \BUS_ADDR_INTERNAL[9]_adj_2 ;
    output \BUS_ADDR_INTERNAL[10]_adj_3 ;
    output \BUS_ADDR_INTERNAL[11]_adj_4 ;
    output \BUS_ADDR_INTERNAL[12]_adj_5 ;
    output \BUS_ADDR_INTERNAL[13]_adj_6 ;
    output \BUS_ADDR_INTERNAL[14]_adj_7 ;
    output \BUS_ADDR_INTERNAL[15]_adj_8 ;
    output \BUS_ADDR_INTERNAL[16]_adj_9 ;
    output \BUS_ADDR_INTERNAL[17] ;
    input PIC_DATA_IN_out_3;
    input PIC_WE_IN_c;
    input PIC_DATA_IN_out_6;
    output n12276;
    output n12274;
    output n12291;
    input \BUS_ADDR_INTERNAL[5]_adj_10 ;
    output n12272;
    input \BUS_ADDR_INTERNAL[6]_adj_11 ;
    output n12289;
    input \BUS_ADDR_INTERNAL[7]_adj_12 ;
    output n12288;
    input PIC_DATA_IN_out_5;
    input PIC_DATA_IN_out_7;
    input \BUS_ADDR_INTERNAL[3]_adj_13 ;
    output n12287;
    output n12290;
    input \BUS_data[4] ;
    input \BUS_data[5] ;
    input \BUS_data[6] ;
    input \BUS_data[7] ;
    input \BUS_ADDR_INTERNAL[1]_adj_14 ;
    output n12292;
    output \writeData[4] ;
    output \writeData[5] ;
    output \writeData[6] ;
    output \writeData[7] ;
    output n12280;
    input n1921;
    output n12222;
    input n2025;
    output LOGIC_CLOCK_enable_26;
    input \BUS_ADDR_INTERNAL[2]_adj_15 ;
    output n12279;
    input \BUS_ADDR_INTERNAL[4]_adj_16 ;
    output n12278;
    input n13147;
    output \state[7] ;
    input \state_7__N_1050[7] ;
    output n12273;
    input n13145;
    input n13146;
    input n13148;
    input n13153;
    input n13149;
    input n13152;
    input \BUS_ADDR_INTERNAL[0]_adj_17 ;
    input n12299;
    input PIC_DATA_IN_out_1;
    input PIC_DATA_IN_out_2;
    input PIC_DATA_IN_out_4;
    output n12223;
    input n13141;
    input n11485;
    input n12219;
    output LOGIC_CLOCK_enable_48;
    output n7167;
    input n12213;
    input n12314;
    output \BUS_DATA_INTERNAL[2] ;
    input n6;
    input \BUS_currGrantID_3__N_72[0] ;
    output \BUS_currGrantID_3__N_72[1] ;
    output n12352;
    output n71;
    input PIC_OE_c;
    output n12312;
    input n12214;
    output n12324;
    input PIC_DATA_IN_out_0;
    input n12212;
    input n12348;
    input n13139;
    output n6_adj_18;
    output \BUS_DATA_INTERNAL[1] ;
    input n10895;
    input n69;
    output n1184;
    output BUS_currGrantID_3__N_54;
    input BUS_DONE;
    output \BUS_DATA_INTERNAL[0] ;
    input n12250;
    input n12217;
    output \PIC_data[9] ;
    output \PIC_data[11] ;
    output \PIC_data[10] ;
    output n100;
    output \PIC_data[12] ;
    output \PIC_data[8] ;
    output \PIC_data[13] ;
    output \PIC_data[14] ;
    input SRAM_WE_N_704;
    input \lastAddress[4] ;
    output n60;
    input n10904;
    input \lastAddress[7] ;
    output n57;
    input \lastAddress[3] ;
    output n61;
    input \lastAddress[17] ;
    output n47;
    input n13140;
    input n12304;
    output lastAddress_31__N_833;
    output lastAddress_31__N_773;
    input n9924;
    output BUS_DONE_OUT_N_626;
    output \BUS_DATA_INTERNAL[3] ;
    input n12332;
    output n10976;
    output n11012;
    
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire BUS_DIRECTION_INTERNAL_N_997 /* synthesis is_clock=1, SET_AS_NETWORK=\PIC_BUS_INTERFACE/BUS_DIRECTION_INTERNAL_N_997 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(38[8:30])
    
    wire n10017;
    wire [7:0]rModDataTrans;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(56[8:21])
    wire [9:0]rModDataWrite_15__N_1120;
    
    wire n10018, n9693;
    wire [18:0]lastAddress;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(41[8:19])
    
    wire n9694, mult_8u_9u_0_cin_lr_0, n10016, n10014;
    wire [16:0]rModDataWrite_15__N_1070;
    wire [15:0]rModDataWrite_15__N_1087;
    wire [16:0]rModDataWrite;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(54[8:21])
    
    wire n12266;
    wire [7:0]state_c;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(48[8:13])
    
    wire n10258, mult_8u_8u_0_cin_lr_0;
    wire [3:0]transferMode;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(50[8:20])
    
    wire LOGIC_CLOCK_enable_116, LOGIC_CLOCK_enable_159;
    wire [7:0]rModDataRead;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(53[8:20])
    
    wire LOGIC_CLOCK_enable_141, BUS_REQ_N_1209;
    wire [15:0]writeData;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(46[8:17])
    
    wire LOGIC_CLOCK_enable_148;
    wire [15:0]writeData_15__N_1169;
    
    wire n10013;
    wire [7:0]state_7__N_1050;
    wire [15:0]data;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(44[8:12])
    
    wire n10012, n11759, n11760, n12233, mult_8u_9u_0_pp_3_16, mult_8u_9u_0_pp_3_15, 
        mco_15, n10011, mult_8u_9u_0_pp_3_14, mult_8u_9u_0_pp_3_13, 
        mco_14, mult_8u_9u_0_pp_3_12, mult_8u_9u_0_pp_3_11, mco_13, 
        mult_8u_9u_0_pp_3_10, mult_8u_9u_0_pp_3_9, mco_12, mult_8u_9u_0_pp_3_8, 
        mult_8u_9u_0_pp_3_7, mult_8u_9u_0_cin_lr_6, n10156, n10155, 
        n4, n14, n23, n10154, n10010, n10153, n10009, n10152, 
        n10008, n10151, n10150, n5334, mult_8u_9u_0_pp_2_14, mult_8u_9u_0_pp_2_13, 
        mco_11, mult_8u_9u_0_pp_2_12, mult_8u_9u_0_pp_2_11, mco_10, 
        mult_8u_9u_0_pp_2_10, mult_8u_9u_0_pp_2_9, mco_9, mult_8u_9u_0_pp_2_8, 
        mult_8u_9u_0_pp_2_7, mco_8, mult_8u_9u_0_pp_2_6, mult_8u_9u_0_pp_2_5, 
        mult_8u_9u_0_cin_lr_4, mult_8u_9u_0_pp_1_12, mult_8u_9u_0_pp_1_11, 
        mco_7, mult_8u_9u_0_pp_1_10, mult_8u_9u_0_pp_1_9, mco_6, mult_8u_9u_0_pp_1_8, 
        mult_8u_9u_0_pp_1_7, mco_5, mult_8u_9u_0_pp_1_6, mult_8u_9u_0_pp_1_5, 
        mco_4, mult_8u_9u_0_pp_1_4, mult_8u_9u_0_pp_1_3, mult_8u_9u_0_cin_lr_2, 
        mult_8u_9u_0_pp_0_10, mult_8u_9u_0_pp_0_9, mco_3, mult_8u_9u_0_pp_0_8, 
        mult_8u_9u_0_pp_0_7, mco_2, mult_8u_9u_0_pp_0_6, mult_8u_9u_0_pp_0_5, 
        mco_1, mult_8u_9u_0_pp_0_4, mult_8u_9u_0_pp_0_3, mco, mult_8u_9u_0_pp_0_2, 
        co_t_mult_8u_9u_0_2_6, s_mult_8u_9u_0_1_15, s_mult_8u_9u_0_1_16, 
        co_t_mult_8u_9u_0_2_5, s_mult_8u_9u_0_1_13, s_mult_8u_9u_0_1_14, 
        s_mult_8u_9u_0_0_13, co_t_mult_8u_9u_0_2_4, s_mult_8u_9u_0_1_11, 
        s_mult_8u_9u_0_1_12, s_mult_8u_9u_0_0_11, s_mult_8u_9u_0_0_12, 
        co_t_mult_8u_9u_0_2_3, s_mult_8u_9u_0_1_9, s_mult_8u_9u_0_1_10, 
        s_mult_8u_9u_0_0_9, s_mult_8u_9u_0_0_10, co_t_mult_8u_9u_0_2_2, 
        s_mult_8u_9u_0_1_7, s_mult_8u_9u_0_1_8, s_mult_8u_9u_0_0_7, s_mult_8u_9u_0_0_8, 
        co_t_mult_8u_9u_0_2_1, s_mult_8u_9u_0_1_6, s_mult_8u_9u_0_0_5, 
        s_mult_8u_9u_0_0_6, mult_8u_9u_0_pp_2_4, s_mult_8u_9u_0_0_4, co_mult_8u_9u_0_1_5, 
        co_mult_8u_9u_0_1_4, co_mult_8u_9u_0_1_3, co_mult_8u_9u_0_1_2, 
        co_mult_8u_9u_0_1_1, mult_8u_9u_0_pp_3_6, co_mult_8u_9u_0_0_6, 
        co_mult_8u_9u_0_0_5, co_mult_8u_9u_0_0_4, co_mult_8u_9u_0_0_3, 
        co_mult_8u_9u_0_0_2, co_mult_8u_9u_0_0_1, mult_8u_9u_0_pp_1_2, 
        LOGIC_CLOCK_enable_46, LOGIC_CLOCK_enable_47, n10891, mult_8u_8u_0_pp_3_6, 
        mult_8u_8u_0_pp_2_4, mult_8u_8u_0_pp_1_2, mult_8u_8u_0_pp_0_9, 
        mfco, mult_8u_8u_0_cin_lr_2, mult_8u_8u_0_pp_1_11, mfco_1, mult_8u_8u_0_cin_lr_4, 
        mult_8u_8u_0_pp_2_13, mfco_2, mult_8u_8u_0_cin_lr_6, mult_8u_8u_0_pp_3_15, 
        mfco_3, co_mult_8u_8u_0_0_1, mult_8u_8u_0_pp_0_2, co_mult_8u_8u_0_0_2, 
        s_mult_8u_8u_0_0_4, mult_8u_8u_0_pp_0_4, mult_8u_8u_0_pp_0_3, 
        mult_8u_8u_0_pp_1_4, mult_8u_8u_0_pp_1_3, co_mult_8u_8u_0_0_3, 
        s_mult_8u_8u_0_0_5, s_mult_8u_8u_0_0_6, mult_8u_8u_0_pp_0_6, mult_8u_8u_0_pp_0_5, 
        mult_8u_8u_0_pp_1_6, mult_8u_8u_0_pp_1_5, co_mult_8u_8u_0_0_4, 
        s_mult_8u_8u_0_0_7, s_mult_8u_8u_0_0_8, mult_8u_8u_0_pp_0_8, mult_8u_8u_0_pp_0_7, 
        mult_8u_8u_0_pp_1_8, mult_8u_8u_0_pp_1_7, co_mult_8u_8u_0_0_5, 
        s_mult_8u_8u_0_0_9, s_mult_8u_8u_0_0_10, mult_8u_8u_0_pp_1_10, 
        mult_8u_8u_0_pp_1_9, co_mult_8u_8u_0_0_6, s_mult_8u_8u_0_0_11, 
        s_mult_8u_8u_0_0_12, s_mult_8u_8u_0_0_13, co_mult_8u_8u_0_1_1, 
        s_mult_8u_8u_0_1_6, mult_8u_8u_0_pp_2_6, co_mult_8u_8u_0_1_2, 
        s_mult_8u_8u_0_1_7, s_mult_8u_8u_0_1_8, mult_8u_8u_0_pp_2_8, mult_8u_8u_0_pp_2_7, 
        mult_8u_8u_0_pp_3_8, mult_8u_8u_0_pp_3_7, co_mult_8u_8u_0_1_3, 
        s_mult_8u_8u_0_1_9, s_mult_8u_8u_0_1_10, mult_8u_8u_0_pp_2_10, 
        mult_8u_8u_0_pp_2_9, mult_8u_8u_0_pp_3_10, mult_8u_8u_0_pp_3_9, 
        co_mult_8u_8u_0_1_4, s_mult_8u_8u_0_1_11, s_mult_8u_8u_0_1_12, 
        mult_8u_8u_0_pp_2_12, mult_8u_8u_0_pp_2_11, mult_8u_8u_0_pp_3_12, 
        mult_8u_8u_0_pp_3_11, co_mult_8u_8u_0_1_5, s_mult_8u_8u_0_1_13, 
        s_mult_8u_8u_0_1_14, mult_8u_8u_0_pp_3_14, mult_8u_8u_0_pp_3_13, 
        s_mult_8u_8u_0_1_15, co_t_mult_8u_8u_0_2_1, co_t_mult_8u_8u_0_2_2, 
        mult_8u_8u_0_pp_2_5, co_t_mult_8u_8u_0_2_3, co_t_mult_8u_8u_0_2_4, 
        co_t_mult_8u_8u_0_2_5, co_t_mult_8u_8u_0_2_6, mco_adj_1242, mco_1_adj_1243, 
        mco_2_adj_1244, mco_3_adj_1245, mco_4_adj_1246, mco_5_adj_1247, 
        mco_6_adj_1248, mco_7_adj_1249, mco_8_adj_1250, mco_9_adj_1251, 
        mco_10_adj_1252, mco_11_adj_1253, n10074, n10073, n10072, 
        n10071, n10070, n10069, n10068, n10067, LOGIC_CLOCK_enable_149, 
        LOGIC_CLOCK_enable_150, LOGIC_CLOCK_enable_151, LOGIC_CLOCK_enable_152, 
        n10066, n10065, n10064, n15, n12236, n12267, n26, n28, 
        n19, n38, n4_adj_1271, n12293, n11014, n11006, n12350, 
        n12351, n11, n12345, BUS_DIRECTION_INTERNAL_N_1000, n11418, 
        n12346, n12323, n12246, n12347, n12245, n12239, n9697, 
        n10324, n23_adj_1273, n16, n10, n8, n12242, n9696, n9695, 
        n10019;
    
    CCU2D add_313_5 (.A0(rModDataTrans[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(rModDataTrans[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10017), .COUT(n10018), .S0(rModDataWrite_15__N_1120[3]), 
          .S1(rModDataWrite_15__N_1120[4]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_313_5.INIT0 = 16'hf555;
    defparam add_313_5.INIT1 = 16'hf555;
    defparam add_313_5.INJECT1_0 = "NO";
    defparam add_313_5.INJECT1_1 = "NO";
    CCU2D lastAddress_18__I_0_13 (.A0(PIC_ADDR_IN_c_15), .B0(lastAddress[15]), 
          .C0(PIC_ADDR_IN_c_14), .D0(lastAddress[14]), .A1(PIC_ADDR_IN_c_13), 
          .B1(lastAddress[13]), .C1(PIC_ADDR_IN_c_12), .D1(lastAddress[12]), 
          .CIN(n9693), .COUT(n9694));
    defparam lastAddress_18__I_0_13.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_13.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_13.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_13.INJECT1_1 = "YES";
    FADD2B mult_8u_9u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    CCU2D add_313_3 (.A0(rModDataTrans[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(rModDataTrans[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10016), .COUT(n10017), .S0(rModDataWrite_15__N_1120[1]), 
          .S1(rModDataWrite_15__N_1120[2]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_313_3.INIT0 = 16'hf555;
    defparam add_313_3.INIT1 = 16'hf555;
    defparam add_313_3.INJECT1_0 = "NO";
    defparam add_313_3.INJECT1_1 = "NO";
    CCU2D add_313_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(rModDataTrans[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n10016), .S1(rModDataWrite_15__N_1120[0]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_313_1.INIT0 = 16'hF000;
    defparam add_313_1.INIT1 = 16'h0aaa;
    defparam add_313_1.INJECT1_0 = "NO";
    defparam add_313_1.INJECT1_1 = "NO";
    CCU2D add_314_16 (.A0(rModDataWrite_15__N_1070[14]), .B0(rModDataWrite_15__N_1087[14]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[15]), 
          .B1(rModDataWrite_15__N_1087[15]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10014), .S0(rModDataWrite[14]), .S1(rModDataWrite[15]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_16.INIT0 = 16'h5666;
    defparam add_314_16.INIT1 = 16'h5666;
    defparam add_314_16.INJECT1_0 = "NO";
    defparam add_314_16.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut (.A(state[1]), .B(n12266), .C(state[4]), .D(state_c[0]), 
         .Z(n10258)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    FADD2B mult_8u_8u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FD1P3AX transferMode_i0_i0 (.D(\BUS_data[0] ), .SP(LOGIC_CLOCK_enable_116), 
            .CK(LOGIC_CLOCK), .Q(transferMode[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i0.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i1 (.D(PIC_ADDR_IN_c_0), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i1.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i0 (.D(\BUS_data[0] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i0.GSR = "DISABLED";
    FD1S3DX BUS_REQ_263 (.D(BUS_REQ_N_1209), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_997), 
            .Q(\BUS_req[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_REQ_263.GSR = "DISABLED";
    FD1P3AX writeData_i0_i0 (.D(writeData_15__N_1169[0]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(writeData[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i0.GSR = "DISABLED";
    CCU2D add_314_14 (.A0(rModDataWrite_15__N_1070[12]), .B0(rModDataWrite_15__N_1087[12]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[13]), 
          .B1(rModDataWrite_15__N_1087[13]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10013), .COUT(n10014), .S0(rModDataWrite[12]), .S1(rModDataWrite[13]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_14.INIT0 = 16'h5666;
    defparam add_314_14.INIT1 = 16'h5666;
    defparam add_314_14.INJECT1_0 = "NO";
    defparam add_314_14.INJECT1_1 = "NO";
    FD1S3DX state_i0 (.D(state_7__N_1050[0]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_997), 
            .Q(state_c[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i0 (.D(data[8]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i0.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i1 (.D(PIC_ADDR_IN_c_0), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i1.GSR = "DISABLED";
    FD1S3DX WRITE_DONE_261 (.D(n13160), .CK(LOGIC_CLOCK), .CD(transferMode_3__N_1115), 
            .Q(WRITE_DONE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam WRITE_DONE_261.GSR = "DISABLED";
    CCU2D add_314_12 (.A0(rModDataWrite_15__N_1070[10]), .B0(rModDataWrite_15__N_1087[10]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[11]), 
          .B1(rModDataWrite_15__N_1087[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10012), .COUT(n10013), .S0(rModDataWrite[10]), .S1(rModDataWrite[11]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_12.INIT0 = 16'h5666;
    defparam add_314_12.INIT1 = 16'h5666;
    defparam add_314_12.INJECT1_0 = "NO";
    defparam add_314_12.INJECT1_1 = "NO";
    FD1S1A PIC_ADDR_IN_18__I_0_i2 (.D(PIC_ADDR_IN_c_1), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i2.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i3 (.D(PIC_ADDR_IN_c_2), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i3.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i4 (.D(PIC_ADDR_IN_c_3), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i4.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i5 (.D(PIC_ADDR_IN_c_4), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i5.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i6 (.D(PIC_ADDR_IN_c_5), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i6.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i7 (.D(PIC_ADDR_IN_c_6), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i7.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i8 (.D(PIC_ADDR_IN_c_7), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i8.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i9 (.D(PIC_ADDR_IN_c_8), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i9.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i10 (.D(PIC_ADDR_IN_c_9), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i10.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i11 (.D(PIC_ADDR_IN_c_10), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i11.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i12 (.D(PIC_ADDR_IN_c_11), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i12.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i13 (.D(PIC_ADDR_IN_c_12), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i13.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i14 (.D(PIC_ADDR_IN_c_13), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i14.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i15 (.D(PIC_ADDR_IN_c_14), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i15.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i16 (.D(PIC_ADDR_IN_c_15), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i16.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i17 (.D(PIC_ADDR_IN_c_16), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[16])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i17.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i18 (.D(PIC_ADDR_IN_c_17), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[17])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i18.GSR = "DISABLED";
    FD1S1A PIC_ADDR_IN_18__I_0_i19 (.D(PIC_ADDR_IN_c_18), .CK(BUS_DIRECTION_INTERNAL_N_997), 
           .Q(lastAddress[18])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(100[2] 157[14])
    defparam PIC_ADDR_IN_18__I_0_i19.GSR = "DISABLED";
    PFUMX i8788 (.BLUT(n11759), .ALUT(n11758), .C0(state[4]), .Z(n11760));
    LUT4 i2_3_lut_4_lut_adj_126 (.A(n12233), .B(n5045), .C(n12252), .D(n12263), 
         .Z(n87)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i2_3_lut_4_lut_adj_126.init = 16'hfeff;
    MULT2 mult_8u_9u_0_mult_6_4 (.A0(rModDataWrite_15__N_1120[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[7]), .B1(rModDataRead[6]), 
          .B2(rModDataRead[7]), .B3(rModDataRead[6]), .CI(mco_15), .P0(mult_8u_9u_0_pp_3_15), 
          .P1(mult_8u_9u_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    CCU2D add_314_10 (.A0(rModDataWrite_15__N_1070[8]), .B0(rModDataWrite_15__N_1087[8]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[9]), 
          .B1(rModDataWrite_15__N_1087[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10011), .COUT(n10012), .S0(rModDataWrite[8]), .S1(rModDataWrite[9]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_10.INIT0 = 16'h5666;
    defparam add_314_10.INIT1 = 16'h5666;
    defparam add_314_10.INJECT1_0 = "NO";
    defparam add_314_10.INJECT1_1 = "NO";
    MULT2 mult_8u_9u_0_mult_6_3 (.A0(rModDataWrite_15__N_1120[6]), .A1(rModDataWrite_15__N_1120[7]), 
          .A2(rModDataWrite_15__N_1120[7]), .A3(rModDataWrite_15__N_1120[8]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mco_14), .CO(mco_15), .P0(mult_8u_9u_0_pp_3_13), 
          .P1(mult_8u_9u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_2 (.A0(rModDataWrite_15__N_1120[4]), .A1(rModDataWrite_15__N_1120[5]), 
          .A2(rModDataWrite_15__N_1120[5]), .A3(rModDataWrite_15__N_1120[6]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mco_13), .CO(mco_14), .P0(mult_8u_9u_0_pp_3_11), 
          .P1(mult_8u_9u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_1 (.A0(rModDataWrite_15__N_1120[2]), .A1(rModDataWrite_15__N_1120[3]), 
          .A2(rModDataWrite_15__N_1120[3]), .A3(rModDataWrite_15__N_1120[4]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mco_12), .CO(mco_13), .P0(mult_8u_9u_0_pp_3_9), 
          .P1(mult_8u_9u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_6_0 (.A0(rModDataWrite_15__N_1120[0]), .A1(rModDataWrite_15__N_1120[1]), 
          .A2(rModDataWrite_15__N_1120[1]), .A3(rModDataWrite_15__N_1120[2]), 
          .B0(rModDataRead[7]), .B1(rModDataRead[6]), .B2(rModDataRead[7]), 
          .B3(rModDataRead[6]), .CI(mult_8u_9u_0_cin_lr_6), .CO(mco_12), 
          .P0(mult_8u_9u_0_pp_3_7), .P1(mult_8u_9u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    CCU2D add_7185_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10156), 
          .S0(BUS_VALID_N_1118));
    defparam add_7185_cout.INIT0 = 16'h0000;
    defparam add_7185_cout.INIT1 = 16'h0000;
    defparam add_7185_cout.INJECT1_0 = "NO";
    defparam add_7185_cout.INJECT1_1 = "NO";
    CCU2D add_7185_13 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n10155), .COUT(n10156));
    defparam add_7185_13.INIT0 = 16'heeee;
    defparam add_7185_13.INIT1 = 16'heeee;
    defparam add_7185_13.INJECT1_0 = "NO";
    defparam add_7185_13.INJECT1_1 = "NO";
    PFUMX i29 (.BLUT(n4), .ALUT(n14), .C0(state_c[0]), .Z(n23));
    CCU2D add_7185_11 (.A0(n13158), .B0(n12344), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), 
          .D1(n12309), .CIN(n10154), .COUT(n10155));
    defparam add_7185_11.INIT0 = 16'h8888;
    defparam add_7185_11.INIT1 = 16'hff20;
    defparam add_7185_11.INJECT1_0 = "NO";
    defparam add_7185_11.INJECT1_1 = "NO";
    CCU2D add_314_8 (.A0(rModDataWrite_15__N_1070[6]), .B0(rModDataWrite_15__N_1087[6]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[7]), 
          .B1(rModDataWrite_15__N_1087[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10010), .COUT(n10011));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_8.INIT0 = 16'h5666;
    defparam add_314_8.INIT1 = 16'h5666;
    defparam add_314_8.INJECT1_0 = "NO";
    defparam add_314_8.INJECT1_1 = "NO";
    CCU2D add_7185_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n13150), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16] ), .D1(n13151), 
          .CIN(n10153), .COUT(n10154));
    defparam add_7185_9.INIT0 = 16'h00ae;
    defparam add_7185_9.INIT1 = 16'h00ae;
    defparam add_7185_9.INJECT1_0 = "NO";
    defparam add_7185_9.INJECT1_1 = "NO";
    CCU2D add_314_6 (.A0(rModDataWrite_15__N_1070[4]), .B0(rModDataWrite_15__N_1087[4]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[5]), 
          .B1(rModDataWrite_15__N_1087[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10009), .COUT(n10010));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_6.INIT0 = 16'h5666;
    defparam add_314_6.INIT1 = 16'h5666;
    defparam add_314_6.INJECT1_0 = "NO";
    defparam add_314_6.INJECT1_1 = "NO";
    CCU2D add_7185_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n13155), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n13157), 
          .CIN(n10152), .COUT(n10153));
    defparam add_7185_7.INIT0 = 16'h00ae;
    defparam add_7185_7.INIT1 = 16'h00ae;
    defparam add_7185_7.INJECT1_0 = "NO";
    defparam add_7185_7.INJECT1_1 = "NO";
    CCU2D add_314_4 (.A0(rModDataWrite_15__N_1070[2]), .B0(rModDataWrite_15__N_1087[2]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[3]), 
          .B1(rModDataWrite_15__N_1087[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n10008), .COUT(n10009));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_4.INIT0 = 16'h5666;
    defparam add_314_4.INIT1 = 16'h5666;
    defparam add_314_4.INJECT1_0 = "NO";
    defparam add_314_4.INJECT1_1 = "NO";
    CCU2D add_7185_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n13156), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n13142), 
          .CIN(n10151), .COUT(n10152));
    defparam add_7185_5.INIT0 = 16'h00ae;
    defparam add_7185_5.INIT1 = 16'h00ae;
    defparam add_7185_5.INJECT1_0 = "NO";
    defparam add_7185_5.INJECT1_1 = "NO";
    CCU2D add_314_2 (.A0(rModDataWrite_15__N_1070[0]), .B0(rModDataWrite_15__N_1087[0]), 
          .C0(GND_net), .D0(GND_net), .A1(rModDataWrite_15__N_1070[1]), 
          .B1(rModDataWrite_15__N_1087[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n10008));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[37:109])
    defparam add_314_2.INIT0 = 16'h7000;
    defparam add_314_2.INIT1 = 16'h5666;
    defparam add_314_2.INJECT1_0 = "NO";
    defparam add_314_2.INJECT1_1 = "NO";
    CCU2D add_7185_3 (.A0(\BUS_ADDR_INTERNAL[9] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13144), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n13143), 
          .CIN(n10150), .COUT(n10151));
    defparam add_7185_3.INIT0 = 16'h00dc;
    defparam add_7185_3.INIT1 = 16'hff51;
    defparam add_7185_3.INJECT1_0 = "NO";
    defparam add_7185_3.INJECT1_1 = "NO";
    CCU2D add_7185_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), 
          .D1(n13154), .COUT(n10150));
    defparam add_7185_1.INIT0 = 16'hF000;
    defparam add_7185_1.INIT1 = 16'h00ae;
    defparam add_7185_1.INJECT1_0 = "NO";
    defparam add_7185_1.INJECT1_1 = "NO";
    FD1P3IX writeData_i0_i15 (.D(PIC_DATA_IN_out_15), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i15.GSR = "DISABLED";
    MULT2 mult_8u_9u_0_mult_4_4 (.A0(rModDataWrite_15__N_1120[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[5]), .B1(rModDataRead[4]), 
          .B2(rModDataRead[5]), .B3(rModDataRead[4]), .CI(mco_11), .P0(mult_8u_9u_0_pp_2_13), 
          .P1(mult_8u_9u_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FD1P3IX writeData_i0_i13 (.D(PIC_DATA_IN_out_13), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i13.GSR = "DISABLED";
    FD1P3IX writeData_i0_i14 (.D(PIC_DATA_IN_out_14), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i14.GSR = "DISABLED";
    MULT2 mult_8u_9u_0_mult_4_3 (.A0(rModDataWrite_15__N_1120[6]), .A1(rModDataWrite_15__N_1120[7]), 
          .A2(rModDataWrite_15__N_1120[7]), .A3(rModDataWrite_15__N_1120[8]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mco_10), .CO(mco_11), .P0(mult_8u_9u_0_pp_2_11), 
          .P1(mult_8u_9u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_2 (.A0(rModDataWrite_15__N_1120[4]), .A1(rModDataWrite_15__N_1120[5]), 
          .A2(rModDataWrite_15__N_1120[5]), .A3(rModDataWrite_15__N_1120[6]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mco_9), .CO(mco_10), .P0(mult_8u_9u_0_pp_2_9), 
          .P1(mult_8u_9u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_1 (.A0(rModDataWrite_15__N_1120[2]), .A1(rModDataWrite_15__N_1120[3]), 
          .A2(rModDataWrite_15__N_1120[3]), .A3(rModDataWrite_15__N_1120[4]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mco_8), .CO(mco_9), .P0(mult_8u_9u_0_pp_2_7), 
          .P1(mult_8u_9u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_4_0 (.A0(rModDataWrite_15__N_1120[0]), .A1(rModDataWrite_15__N_1120[1]), 
          .A2(rModDataWrite_15__N_1120[1]), .A3(rModDataWrite_15__N_1120[2]), 
          .B0(rModDataRead[5]), .B1(rModDataRead[4]), .B2(rModDataRead[5]), 
          .B3(rModDataRead[4]), .CI(mult_8u_9u_0_cin_lr_4), .CO(mco_8), 
          .P0(mult_8u_9u_0_pp_2_5), .P1(mult_8u_9u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_4 (.A0(rModDataWrite_15__N_1120[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[3]), .B1(rModDataRead[2]), 
          .B2(rModDataRead[3]), .B3(rModDataRead[2]), .CI(mco_7), .P0(mult_8u_9u_0_pp_1_11), 
          .P1(mult_8u_9u_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_3 (.A0(rModDataWrite_15__N_1120[6]), .A1(rModDataWrite_15__N_1120[7]), 
          .A2(rModDataWrite_15__N_1120[7]), .A3(rModDataWrite_15__N_1120[8]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mco_6), .CO(mco_7), .P0(mult_8u_9u_0_pp_1_9), 
          .P1(mult_8u_9u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FD1P3IX writeData_i0_i11 (.D(PIC_DATA_IN_out_11), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i11.GSR = "DISABLED";
    FD1P3IX writeData_i0_i12 (.D(PIC_DATA_IN_out_12), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i12.GSR = "DISABLED";
    MULT2 mult_8u_9u_0_mult_2_2 (.A0(rModDataWrite_15__N_1120[4]), .A1(rModDataWrite_15__N_1120[5]), 
          .A2(rModDataWrite_15__N_1120[5]), .A3(rModDataWrite_15__N_1120[6]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mco_5), .CO(mco_6), .P0(mult_8u_9u_0_pp_1_7), 
          .P1(mult_8u_9u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_1 (.A0(rModDataWrite_15__N_1120[2]), .A1(rModDataWrite_15__N_1120[3]), 
          .A2(rModDataWrite_15__N_1120[3]), .A3(rModDataWrite_15__N_1120[4]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mco_4), .CO(mco_5), .P0(mult_8u_9u_0_pp_1_5), 
          .P1(mult_8u_9u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_2_0 (.A0(rModDataWrite_15__N_1120[0]), .A1(rModDataWrite_15__N_1120[1]), 
          .A2(rModDataWrite_15__N_1120[1]), .A3(rModDataWrite_15__N_1120[2]), 
          .B0(rModDataRead[3]), .B1(rModDataRead[2]), .B2(rModDataRead[3]), 
          .B3(rModDataRead[2]), .CI(mult_8u_9u_0_cin_lr_2), .CO(mco_4), 
          .P0(mult_8u_9u_0_pp_1_3), .P1(mult_8u_9u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_4 (.A0(rModDataWrite_15__N_1120[8]), .A1(GND_net), 
          .A2(GND_net), .A3(GND_net), .B0(rModDataRead[1]), .B1(rModDataRead[0]), 
          .B2(rModDataRead[1]), .B3(rModDataRead[0]), .CI(mco_3), .P0(mult_8u_9u_0_pp_0_9), 
          .P1(mult_8u_9u_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_3 (.A0(rModDataWrite_15__N_1120[6]), .A1(rModDataWrite_15__N_1120[7]), 
          .A2(rModDataWrite_15__N_1120[7]), .A3(rModDataWrite_15__N_1120[8]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mco_2), .CO(mco_3), .P0(mult_8u_9u_0_pp_0_7), 
          .P1(mult_8u_9u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_2 (.A0(rModDataWrite_15__N_1120[4]), .A1(rModDataWrite_15__N_1120[5]), 
          .A2(rModDataWrite_15__N_1120[5]), .A3(rModDataWrite_15__N_1120[6]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mco_1), .CO(mco_2), .P0(mult_8u_9u_0_pp_0_5), 
          .P1(mult_8u_9u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FD1P3IX writeData_i0_i9 (.D(PIC_DATA_IN_out_9), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i9.GSR = "DISABLED";
    FD1P3IX writeData_i0_i10 (.D(PIC_DATA_IN_out_10), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i10.GSR = "DISABLED";
    MULT2 mult_8u_9u_0_mult_0_1 (.A0(rModDataWrite_15__N_1120[2]), .A1(rModDataWrite_15__N_1120[3]), 
          .A2(rModDataWrite_15__N_1120[3]), .A3(rModDataWrite_15__N_1120[4]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mco), .CO(mco_1), .P0(mult_8u_9u_0_pp_0_3), 
          .P1(mult_8u_9u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    MULT2 mult_8u_9u_0_mult_0_0 (.A0(rModDataWrite_15__N_1120[0]), .A1(rModDataWrite_15__N_1120[1]), 
          .A2(rModDataWrite_15__N_1120[1]), .A3(rModDataWrite_15__N_1120[2]), 
          .B0(rModDataRead[1]), .B1(rModDataRead[0]), .B2(rModDataRead[1]), 
          .B3(rModDataRead[0]), .CI(mult_8u_9u_0_cin_lr_0), .CO(mco), 
          .P0(rModDataWrite_15__N_1070[1]), .P1(mult_8u_9u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_7 (.A0(GND_net), .A1(GND_net), .B0(s_mult_8u_9u_0_1_15), 
           .B1(s_mult_8u_9u_0_1_16), .CI(co_t_mult_8u_9u_0_2_6), .S0(rModDataWrite_15__N_1070[15])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_6 (.A0(s_mult_8u_9u_0_0_13), .A1(GND_net), 
           .B0(s_mult_8u_9u_0_1_13), .B1(s_mult_8u_9u_0_1_14), .CI(co_t_mult_8u_9u_0_2_5), 
           .COUT(co_t_mult_8u_9u_0_2_6), .S0(rModDataWrite_15__N_1070[13]), 
           .S1(rModDataWrite_15__N_1070[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_5 (.A0(s_mult_8u_9u_0_0_11), .A1(s_mult_8u_9u_0_0_12), 
           .B0(s_mult_8u_9u_0_1_11), .B1(s_mult_8u_9u_0_1_12), .CI(co_t_mult_8u_9u_0_2_4), 
           .COUT(co_t_mult_8u_9u_0_2_5), .S0(rModDataWrite_15__N_1070[11]), 
           .S1(rModDataWrite_15__N_1070[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FD1P3IX writeData_i0_i8 (.D(PIC_DATA_IN_out_8), .SP(LOGIC_CLOCK_enable_148), 
            .CD(n5334), .CK(LOGIC_CLOCK), .Q(writeData[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i8.GSR = "DISABLED";
    FADD2B t_mult_8u_9u_0_add_2_4 (.A0(s_mult_8u_9u_0_0_9), .A1(s_mult_8u_9u_0_0_10), 
           .B0(s_mult_8u_9u_0_1_9), .B1(s_mult_8u_9u_0_1_10), .CI(co_t_mult_8u_9u_0_2_3), 
           .COUT(co_t_mult_8u_9u_0_2_4), .S0(rModDataWrite_15__N_1070[9]), 
           .S1(rModDataWrite_15__N_1070[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_3 (.A0(s_mult_8u_9u_0_0_7), .A1(s_mult_8u_9u_0_0_8), 
           .B0(s_mult_8u_9u_0_1_7), .B1(s_mult_8u_9u_0_1_8), .CI(co_t_mult_8u_9u_0_2_2), 
           .COUT(co_t_mult_8u_9u_0_2_3), .S0(rModDataWrite_15__N_1070[7]), 
           .S1(rModDataWrite_15__N_1070[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B t_mult_8u_9u_0_add_2_2 (.A0(s_mult_8u_9u_0_0_5), .A1(s_mult_8u_9u_0_0_6), 
           .B0(mult_8u_9u_0_pp_2_5), .B1(s_mult_8u_9u_0_1_6), .CI(co_t_mult_8u_9u_0_2_1), 
           .COUT(co_t_mult_8u_9u_0_2_2), .S0(rModDataWrite_15__N_1070[5]), 
           .S1(rModDataWrite_15__N_1070[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_t_mult_8u_9u_0_2_1 (.A0(GND_net), .A1(s_mult_8u_9u_0_0_4), 
           .B0(GND_net), .B1(mult_8u_9u_0_pp_2_4), .CI(GND_net), .COUT(co_t_mult_8u_9u_0_2_1), 
           .S1(rModDataWrite_15__N_1070[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_9u_0_pp_3_15), 
           .B1(mult_8u_9u_0_pp_3_16), .CI(co_mult_8u_9u_0_1_5), .S0(s_mult_8u_9u_0_1_15), 
           .S1(s_mult_8u_9u_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_5 (.A0(mult_8u_9u_0_pp_2_13), .A1(mult_8u_9u_0_pp_2_14), 
           .B0(mult_8u_9u_0_pp_3_13), .B1(mult_8u_9u_0_pp_3_14), .CI(co_mult_8u_9u_0_1_4), 
           .COUT(co_mult_8u_9u_0_1_5), .S0(s_mult_8u_9u_0_1_13), .S1(s_mult_8u_9u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_4 (.A0(mult_8u_9u_0_pp_2_11), .A1(mult_8u_9u_0_pp_2_12), 
           .B0(mult_8u_9u_0_pp_3_11), .B1(mult_8u_9u_0_pp_3_12), .CI(co_mult_8u_9u_0_1_3), 
           .COUT(co_mult_8u_9u_0_1_4), .S0(s_mult_8u_9u_0_1_11), .S1(s_mult_8u_9u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_3 (.A0(mult_8u_9u_0_pp_2_9), .A1(mult_8u_9u_0_pp_2_10), 
           .B0(mult_8u_9u_0_pp_3_9), .B1(mult_8u_9u_0_pp_3_10), .CI(co_mult_8u_9u_0_1_2), 
           .COUT(co_mult_8u_9u_0_1_3), .S0(s_mult_8u_9u_0_1_9), .S1(s_mult_8u_9u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_1_2 (.A0(mult_8u_9u_0_pp_2_7), .A1(mult_8u_9u_0_pp_2_8), 
           .B0(mult_8u_9u_0_pp_3_7), .B1(mult_8u_9u_0_pp_3_8), .CI(co_mult_8u_9u_0_1_1), 
           .COUT(co_mult_8u_9u_0_1_2), .S0(s_mult_8u_9u_0_1_7), .S1(s_mult_8u_9u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_mult_8u_9u_0_1_1 (.A0(GND_net), .A1(mult_8u_9u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_8u_9u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_8u_9u_0_1_1), 
           .S1(s_mult_8u_9u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_mult_8u_9u_0_0_7 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_8u_9u_0_0_6), .S0(s_mult_8u_9u_0_0_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_9u_0_pp_1_11), 
           .B1(mult_8u_9u_0_pp_1_12), .CI(co_mult_8u_9u_0_0_5), .COUT(co_mult_8u_9u_0_0_6), 
           .S0(s_mult_8u_9u_0_0_11), .S1(s_mult_8u_9u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    CCU2D lastAddress_18__I_0_0 (.A0(PIC_ADDR_IN_c_18), .B0(lastAddress[18]), 
          .C0(GND_net), .D0(GND_net), .A1(PIC_ADDR_IN_c_17), .B1(lastAddress[17]), 
          .C1(PIC_ADDR_IN_c_16), .D1(lastAddress[16]), .COUT(n9693));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[57:82])
    defparam lastAddress_18__I_0_0.INIT0 = 16'h9000;
    defparam lastAddress_18__I_0_0.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_0.INJECT1_0 = "NO";
    defparam lastAddress_18__I_0_0.INJECT1_1 = "YES";
    FADD2B mult_8u_9u_0_add_0_5 (.A0(mult_8u_9u_0_pp_0_9), .A1(mult_8u_9u_0_pp_0_10), 
           .B0(mult_8u_9u_0_pp_1_9), .B1(mult_8u_9u_0_pp_1_10), .CI(co_mult_8u_9u_0_0_4), 
           .COUT(co_mult_8u_9u_0_0_5), .S0(s_mult_8u_9u_0_0_9), .S1(s_mult_8u_9u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_4 (.A0(mult_8u_9u_0_pp_0_7), .A1(mult_8u_9u_0_pp_0_8), 
           .B0(mult_8u_9u_0_pp_1_7), .B1(mult_8u_9u_0_pp_1_8), .CI(co_mult_8u_9u_0_0_3), 
           .COUT(co_mult_8u_9u_0_0_4), .S0(s_mult_8u_9u_0_0_7), .S1(s_mult_8u_9u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_3 (.A0(mult_8u_9u_0_pp_0_5), .A1(mult_8u_9u_0_pp_0_6), 
           .B0(mult_8u_9u_0_pp_1_5), .B1(mult_8u_9u_0_pp_1_6), .CI(co_mult_8u_9u_0_0_2), 
           .COUT(co_mult_8u_9u_0_0_3), .S0(s_mult_8u_9u_0_0_5), .S1(s_mult_8u_9u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_add_0_2 (.A0(mult_8u_9u_0_pp_0_3), .A1(mult_8u_9u_0_pp_0_4), 
           .B0(mult_8u_9u_0_pp_1_3), .B1(mult_8u_9u_0_pp_1_4), .CI(co_mult_8u_9u_0_0_1), 
           .COUT(co_mult_8u_9u_0_0_2), .S0(rModDataWrite_15__N_1070[3]), 
           .S1(s_mult_8u_9u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B Cadd_mult_8u_9u_0_0_1 (.A0(GND_net), .A1(mult_8u_9u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_8u_9u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_8u_9u_0_0_1), 
           .S1(rModDataWrite_15__N_1070[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FADD2B mult_8u_9u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_9u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:108])
    FD1P3DX PIC_READY_264 (.D(n13160), .SP(LOGIC_CLOCK_enable_46), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_997), .Q(PIC_READY_c)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam PIC_READY_264.GSR = "DISABLED";
    AND2 AND2_t3 (.A(rModDataWrite_15__N_1120[0]), .B(rModDataRead[0]), 
         .Z(rModDataWrite_15__N_1070[0])) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(128[10:63])
    AND2 AND2_t2 (.A(rModDataWrite_15__N_1120[0]), .B(rModDataRead[2]), 
         .Z(mult_8u_9u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(130[10:63])
    AND2 AND2_t1 (.A(rModDataWrite_15__N_1120[0]), .B(rModDataRead[4]), 
         .Z(mult_8u_9u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(132[10:63])
    AND2 AND2_t0 (.A(rModDataWrite_15__N_1120[0]), .B(rModDataRead[6]), 
         .Z(mult_8u_9u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_9u.v(134[10:63])
    FD1P3AX BUS_DIRECTION_INTERNAL_269 (.D(n10891), .SP(LOGIC_CLOCK_enable_47), 
            .CK(LOGIC_CLOCK), .Q(BUS_DIRECTION_INTERNAL)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_DIRECTION_INTERNAL_269.GSR = "DISABLED";
    AND2 AND2_t0_adj_127 (.A(data[0]), .B(rModDataTrans[6]), .Z(mult_8u_8u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(125[10:63])
    AND2 AND2_t1_adj_128 (.A(data[0]), .B(rModDataTrans[4]), .Z(mult_8u_8u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(123[10:63])
    AND2 AND2_t2_adj_129 (.A(data[0]), .B(rModDataTrans[2]), .Z(mult_8u_8u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(121[10:63])
    AND2 AND2_t3_adj_130 (.A(data[0]), .B(rModDataTrans[0]), .Z(rModDataWrite_15__N_1087[0])) /* synthesis syn_instantiated=1 */ ;   // mult_8u_8u.v(119[10:63])
    FADD2B mult_8u_8u_0_Cadd_0_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco), .S0(mult_8u_8u_0_pp_0_9)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_Cadd_2_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_1), .S0(mult_8u_8u_0_pp_1_11)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_Cadd_4_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_2), .S0(mult_8u_8u_0_pp_2_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_8u_8u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_Cadd_6_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(mfco_3), .S0(mult_8u_8u_0_pp_3_15)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_mult_8u_8u_0_0_1 (.A0(GND_net), .A1(mult_8u_8u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_8u_8u_0_0_1), 
           .S1(rModDataWrite_15__N_1087[2])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_2 (.A0(mult_8u_8u_0_pp_0_3), .A1(mult_8u_8u_0_pp_0_4), 
           .B0(mult_8u_8u_0_pp_1_3), .B1(mult_8u_8u_0_pp_1_4), .CI(co_mult_8u_8u_0_0_1), 
           .COUT(co_mult_8u_8u_0_0_2), .S0(rModDataWrite_15__N_1087[3]), 
           .S1(s_mult_8u_8u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_3 (.A0(mult_8u_8u_0_pp_0_5), .A1(mult_8u_8u_0_pp_0_6), 
           .B0(mult_8u_8u_0_pp_1_5), .B1(mult_8u_8u_0_pp_1_6), .CI(co_mult_8u_8u_0_0_2), 
           .COUT(co_mult_8u_8u_0_0_3), .S0(s_mult_8u_8u_0_0_5), .S1(s_mult_8u_8u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_4 (.A0(mult_8u_8u_0_pp_0_7), .A1(mult_8u_8u_0_pp_0_8), 
           .B0(mult_8u_8u_0_pp_1_7), .B1(mult_8u_8u_0_pp_1_8), .CI(co_mult_8u_8u_0_0_3), 
           .COUT(co_mult_8u_8u_0_0_4), .S0(s_mult_8u_8u_0_0_7), .S1(s_mult_8u_8u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_5 (.A0(mult_8u_8u_0_pp_0_9), .A1(GND_net), 
           .B0(mult_8u_8u_0_pp_1_9), .B1(mult_8u_8u_0_pp_1_10), .CI(co_mult_8u_8u_0_0_4), 
           .COUT(co_mult_8u_8u_0_0_5), .S0(s_mult_8u_8u_0_0_9), .S1(s_mult_8u_8u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_0_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_8u_0_pp_1_11), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_0_5), .COUT(co_mult_8u_8u_0_0_6), 
           .S0(s_mult_8u_8u_0_0_11), .S1(s_mult_8u_8u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_mult_8u_8u_0_0_7 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_0_6), .S0(s_mult_8u_8u_0_0_13)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_mult_8u_8u_0_1_1 (.A0(GND_net), .A1(mult_8u_8u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_8u_8u_0_1_1), 
           .S1(s_mult_8u_8u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_2 (.A0(mult_8u_8u_0_pp_2_7), .A1(mult_8u_8u_0_pp_2_8), 
           .B0(mult_8u_8u_0_pp_3_7), .B1(mult_8u_8u_0_pp_3_8), .CI(co_mult_8u_8u_0_1_1), 
           .COUT(co_mult_8u_8u_0_1_2), .S0(s_mult_8u_8u_0_1_7), .S1(s_mult_8u_8u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_3 (.A0(mult_8u_8u_0_pp_2_9), .A1(mult_8u_8u_0_pp_2_10), 
           .B0(mult_8u_8u_0_pp_3_9), .B1(mult_8u_8u_0_pp_3_10), .CI(co_mult_8u_8u_0_1_2), 
           .COUT(co_mult_8u_8u_0_1_3), .S0(s_mult_8u_8u_0_1_9), .S1(s_mult_8u_8u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_4 (.A0(mult_8u_8u_0_pp_2_11), .A1(mult_8u_8u_0_pp_2_12), 
           .B0(mult_8u_8u_0_pp_3_11), .B1(mult_8u_8u_0_pp_3_12), .CI(co_mult_8u_8u_0_1_3), 
           .COUT(co_mult_8u_8u_0_1_4), .S0(s_mult_8u_8u_0_1_11), .S1(s_mult_8u_8u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_5 (.A0(mult_8u_8u_0_pp_2_13), .A1(GND_net), 
           .B0(mult_8u_8u_0_pp_3_13), .B1(mult_8u_8u_0_pp_3_14), .CI(co_mult_8u_8u_0_1_4), 
           .COUT(co_mult_8u_8u_0_1_5), .S0(s_mult_8u_8u_0_1_13), .S1(s_mult_8u_8u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B mult_8u_8u_0_add_1_6 (.A0(GND_net), .A1(GND_net), .B0(mult_8u_8u_0_pp_3_15), 
           .B1(GND_net), .CI(co_mult_8u_8u_0_1_5), .S0(s_mult_8u_8u_0_1_15)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B Cadd_t_mult_8u_8u_0_2_1 (.A0(GND_net), .A1(s_mult_8u_8u_0_0_4), 
           .B0(GND_net), .B1(mult_8u_8u_0_pp_2_4), .CI(GND_net), .COUT(co_t_mult_8u_8u_0_2_1), 
           .S1(rModDataWrite_15__N_1087[4])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_2 (.A0(s_mult_8u_8u_0_0_5), .A1(s_mult_8u_8u_0_0_6), 
           .B0(mult_8u_8u_0_pp_2_5), .B1(s_mult_8u_8u_0_1_6), .CI(co_t_mult_8u_8u_0_2_1), 
           .COUT(co_t_mult_8u_8u_0_2_2), .S0(rModDataWrite_15__N_1087[5]), 
           .S1(rModDataWrite_15__N_1087[6])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_3 (.A0(s_mult_8u_8u_0_0_7), .A1(s_mult_8u_8u_0_0_8), 
           .B0(s_mult_8u_8u_0_1_7), .B1(s_mult_8u_8u_0_1_8), .CI(co_t_mult_8u_8u_0_2_2), 
           .COUT(co_t_mult_8u_8u_0_2_3), .S0(rModDataWrite_15__N_1087[7]), 
           .S1(rModDataWrite_15__N_1087[8])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_4 (.A0(s_mult_8u_8u_0_0_9), .A1(s_mult_8u_8u_0_0_10), 
           .B0(s_mult_8u_8u_0_1_9), .B1(s_mult_8u_8u_0_1_10), .CI(co_t_mult_8u_8u_0_2_3), 
           .COUT(co_t_mult_8u_8u_0_2_4), .S0(rModDataWrite_15__N_1087[9]), 
           .S1(rModDataWrite_15__N_1087[10])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_5 (.A0(s_mult_8u_8u_0_0_11), .A1(s_mult_8u_8u_0_0_12), 
           .B0(s_mult_8u_8u_0_1_11), .B1(s_mult_8u_8u_0_1_12), .CI(co_t_mult_8u_8u_0_2_4), 
           .COUT(co_t_mult_8u_8u_0_2_5), .S0(rModDataWrite_15__N_1087[11]), 
           .S1(rModDataWrite_15__N_1087[12])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_6 (.A0(s_mult_8u_8u_0_0_13), .A1(GND_net), 
           .B0(s_mult_8u_8u_0_1_13), .B1(s_mult_8u_8u_0_1_14), .CI(co_t_mult_8u_8u_0_2_5), 
           .COUT(co_t_mult_8u_8u_0_2_6), .S0(rModDataWrite_15__N_1087[13]), 
           .S1(rModDataWrite_15__N_1087[14])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    FADD2B t_mult_8u_8u_0_add_2_7 (.A0(GND_net), .A1(GND_net), .B0(s_mult_8u_8u_0_1_15), 
           .B1(GND_net), .CI(co_t_mult_8u_8u_0_2_6), .S0(rModDataWrite_15__N_1087[15])) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_0 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mult_8u_8u_0_cin_lr_0), 
          .CO(mco_adj_1242), .P0(rModDataWrite_15__N_1087[1]), .P1(mult_8u_8u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_1 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mco_adj_1242), 
          .CO(mco_1_adj_1243), .P0(mult_8u_8u_0_pp_0_3), .P1(mult_8u_8u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_2 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mco_1_adj_1243), 
          .CO(mco_2_adj_1244), .P0(mult_8u_8u_0_pp_0_5), .P1(mult_8u_8u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_0_3 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[1]), .B1(rModDataTrans[0]), 
          .B2(rModDataTrans[1]), .B3(rModDataTrans[0]), .CI(mco_2_adj_1244), 
          .CO(mfco), .P0(mult_8u_8u_0_pp_0_7), .P1(mult_8u_8u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_0 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mult_8u_8u_0_cin_lr_2), 
          .CO(mco_3_adj_1245), .P0(mult_8u_8u_0_pp_1_3), .P1(mult_8u_8u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_1 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mco_3_adj_1245), 
          .CO(mco_4_adj_1246), .P0(mult_8u_8u_0_pp_1_5), .P1(mult_8u_8u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_2 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mco_4_adj_1246), 
          .CO(mco_5_adj_1247), .P0(mult_8u_8u_0_pp_1_7), .P1(mult_8u_8u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_2_3 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[3]), .B1(rModDataTrans[2]), 
          .B2(rModDataTrans[3]), .B3(rModDataTrans[2]), .CI(mco_5_adj_1247), 
          .CO(mfco_1), .P0(mult_8u_8u_0_pp_1_9), .P1(mult_8u_8u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_0 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mult_8u_8u_0_cin_lr_4), 
          .CO(mco_6_adj_1248), .P0(mult_8u_8u_0_pp_2_5), .P1(mult_8u_8u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_1 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mco_6_adj_1248), 
          .CO(mco_7_adj_1249), .P0(mult_8u_8u_0_pp_2_7), .P1(mult_8u_8u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_2 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mco_7_adj_1249), 
          .CO(mco_8_adj_1250), .P0(mult_8u_8u_0_pp_2_9), .P1(mult_8u_8u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_4_3 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[5]), .B1(rModDataTrans[4]), 
          .B2(rModDataTrans[5]), .B3(rModDataTrans[4]), .CI(mco_8_adj_1250), 
          .CO(mfco_2), .P0(mult_8u_8u_0_pp_2_11), .P1(mult_8u_8u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_0 (.A0(data[0]), .A1(data[1]), .A2(data[1]), 
          .A3(data[2]), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mult_8u_8u_0_cin_lr_6), 
          .CO(mco_9_adj_1251), .P0(mult_8u_8u_0_pp_3_7), .P1(mult_8u_8u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_1 (.A0(data[2]), .A1(data[3]), .A2(data[3]), 
          .A3(data[4]), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mco_9_adj_1251), 
          .CO(mco_10_adj_1252), .P0(mult_8u_8u_0_pp_3_9), .P1(mult_8u_8u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_2 (.A0(data[4]), .A1(data[5]), .A2(data[5]), 
          .A3(data[6]), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mco_10_adj_1252), 
          .CO(mco_11_adj_1253), .P0(mult_8u_8u_0_pp_3_11), .P1(mult_8u_8u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    MULT2 mult_8u_8u_0_mult_6_3 (.A0(data[6]), .A1(data[7]), .A2(data[7]), 
          .A3(GND_net), .B0(rModDataTrans[7]), .B1(rModDataTrans[6]), 
          .B2(rModDataTrans[7]), .B3(rModDataTrans[6]), .CI(mco_11_adj_1253), 
          .CO(mfco_3), .P0(mult_8u_8u_0_pp_3_13), .P1(mult_8u_8u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[143:166])
    CCU2D add_7189_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10074), 
          .S0(n2198));
    defparam add_7189_cout.INIT0 = 16'h0000;
    defparam add_7189_cout.INIT1 = 16'h0000;
    defparam add_7189_cout.INJECT1_0 = "NO";
    defparam add_7189_cout.INJECT1_1 = "NO";
    FD1P3AX transferMode_i0_i1 (.D(\BUS_data[1] ), .SP(LOGIC_CLOCK_enable_116), 
            .CK(LOGIC_CLOCK), .Q(transferMode[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i1.GSR = "DISABLED";
    FD1P3AX transferMode_i0_i2 (.D(\BUS_data[2] ), .SP(LOGIC_CLOCK_enable_116), 
            .CK(LOGIC_CLOCK), .Q(transferMode[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i2.GSR = "DISABLED";
    FD1P3AX transferMode_i0_i3 (.D(\BUS_data[3] ), .SP(LOGIC_CLOCK_enable_116), 
            .CK(LOGIC_CLOCK), .Q(transferMode[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(80[3] 87[10])
    defparam transferMode_i0_i3.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i2 (.D(PIC_ADDR_IN_c_1), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i2.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i3 (.D(PIC_ADDR_IN_c_2), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i3.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i4 (.D(PIC_ADDR_IN_c_3), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i4.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i5 (.D(PIC_ADDR_IN_c_4), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i5.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i6 (.D(PIC_ADDR_IN_c_5), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i6.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i7 (.D(PIC_ADDR_IN_c_6), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i7.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i8 (.D(PIC_ADDR_IN_c_7), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i8.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i9 (.D(PIC_ADDR_IN_c_8), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[8]_adj_1 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i9.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i10 (.D(PIC_ADDR_IN_c_9), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[9]_adj_2 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i10.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i11 (.D(PIC_ADDR_IN_c_10), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[10]_adj_3 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i11.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i12 (.D(PIC_ADDR_IN_c_11), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[11]_adj_4 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i12.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i13 (.D(PIC_ADDR_IN_c_12), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[12]_adj_5 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i13.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i14 (.D(PIC_ADDR_IN_c_13), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[13]_adj_6 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i14.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i15 (.D(PIC_ADDR_IN_c_14), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[14]_adj_7 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i15.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i16 (.D(PIC_ADDR_IN_c_15), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[15]_adj_8 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i16.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i17 (.D(PIC_ADDR_IN_c_16), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[16]_adj_9 )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i17.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i18 (.D(PIC_ADDR_IN_c_17), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i18.GSR = "DISABLED";
    FD1P3AX BUS_ADDR_INTERNAL__i19 (.D(PIC_ADDR_IN_c_18), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(\BUS_ADDR_INTERNAL[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam BUS_ADDR_INTERNAL__i19.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i1 (.D(\BUS_data[1] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i1.GSR = "DISABLED";
    CCU2D add_7189_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n10073), .COUT(n10074));
    defparam add_7189_21.INIT0 = 16'heeee;
    defparam add_7189_21.INIT1 = 16'heeee;
    defparam add_7189_21.INJECT1_0 = "NO";
    defparam add_7189_21.INJECT1_1 = "NO";
    LUT4 i4809_2_lut (.A(PIC_DATA_IN_out_3), .B(PIC_WE_IN_c), .Z(data[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4809_2_lut.init = 16'h2222;
    LUT4 i4812_2_lut (.A(PIC_DATA_IN_out_6), .B(PIC_WE_IN_c), .Z(data[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4812_2_lut.init = 16'h2222;
    LUT4 PIC_addr_31__I_0_i13_3_lut_rep_250_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[12]_adj_5 ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[12] ), 
         .Z(n12276)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam PIC_addr_31__I_0_i13_3_lut_rep_250_4_lut_4_lut.init = 16'h3808;
    LUT4 i1_3_lut_rep_248_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[10]_adj_3 ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[10] ), 
         .Z(n12274)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_248_4_lut_4_lut.init = 16'h3808;
    LUT4 i1_3_lut_rep_265_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[9]_adj_2 ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[9] ), .Z(n12291)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_265_4_lut_4_lut.init = 16'h3808;
    LUT4 i1_3_lut_rep_246_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[5] ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[5]_adj_10 ), .Z(n12272)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_246_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i7_3_lut_rep_263_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[6] ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[6]_adj_11 ), 
         .Z(n12289)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam PIC_addr_31__I_0_i7_3_lut_rep_263_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i8_3_lut_rep_262_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[7] ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[7]_adj_12 ), 
         .Z(n12288)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam PIC_addr_31__I_0_i8_3_lut_rep_262_4_lut_4_lut.init = 16'h3808;
    LUT4 i4811_2_lut (.A(PIC_DATA_IN_out_5), .B(PIC_WE_IN_c), .Z(data[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4811_2_lut.init = 16'h2222;
    LUT4 i4813_2_lut (.A(PIC_DATA_IN_out_7), .B(PIC_WE_IN_c), .Z(data[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4813_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_rep_261_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[3] ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[3]_adj_13 ), .Z(n12287)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_261_4_lut_4_lut.init = 16'h3808;
    LUT4 PIC_addr_31__I_0_i16_3_lut_rep_264_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[15]_adj_8 ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[15] ), 
         .Z(n12290)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam PIC_addr_31__I_0_i16_3_lut_rep_264_4_lut_4_lut.init = 16'h3808;
    CCU2D add_7189_19 (.A0(n13158), .B0(n12344), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), 
          .D1(n12309), .CIN(n10072), .COUT(n10073));
    defparam add_7189_19.INIT0 = 16'h8888;
    defparam add_7189_19.INIT1 = 16'hff20;
    defparam add_7189_19.INJECT1_0 = "NO";
    defparam add_7189_19.INJECT1_1 = "NO";
    CCU2D add_7189_17 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n13150), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16] ), .D1(n13151), 
          .CIN(n10071), .COUT(n10072));
    defparam add_7189_17.INIT0 = 16'h00ae;
    defparam add_7189_17.INIT1 = 16'h00ae;
    defparam add_7189_17.INJECT1_0 = "NO";
    defparam add_7189_17.INJECT1_1 = "NO";
    CCU2D add_7189_15 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n13155), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n13157), 
          .CIN(n10070), .COUT(n10071));
    defparam add_7189_15.INIT0 = 16'h00ae;
    defparam add_7189_15.INIT1 = 16'h00ae;
    defparam add_7189_15.INJECT1_0 = "NO";
    defparam add_7189_15.INJECT1_1 = "NO";
    FD1P3AX rModDataRead_i0_i2 (.D(\BUS_data[2] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i2.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i3 (.D(\BUS_data[3] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i3.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i4 (.D(\BUS_data[4] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i4.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i5 (.D(\BUS_data[5] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i5.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i6 (.D(\BUS_data[6] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i6.GSR = "DISABLED";
    FD1P3AX rModDataRead_i0_i7 (.D(\BUS_data[7] ), .SP(LOGIC_CLOCK_enable_141), 
            .CK(LOGIC_CLOCK), .Q(rModDataRead[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataRead_i0_i7.GSR = "DISABLED";
    FD1P3AX writeData_i0_i1 (.D(writeData_15__N_1169[1]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(writeData[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i1.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_266_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[1] ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[1]_adj_14 ), .Z(n12292)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_266_4_lut_4_lut.init = 16'h3808;
    FD1P3AX writeData_i0_i2 (.D(writeData_15__N_1169[2]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(writeData[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i2.GSR = "DISABLED";
    FD1P3AX writeData_i0_i3 (.D(writeData_15__N_1169[3]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(writeData[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i3.GSR = "DISABLED";
    FD1P3AX writeData_i0_i4 (.D(writeData_15__N_1169[4]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(\writeData[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i4.GSR = "DISABLED";
    FD1P3AX writeData_i0_i5 (.D(writeData_15__N_1169[5]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(\writeData[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i5.GSR = "DISABLED";
    FD1P3AX writeData_i0_i6 (.D(writeData_15__N_1169[6]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(\writeData[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i6.GSR = "DISABLED";
    FD1P3AX writeData_i0_i7 (.D(writeData_15__N_1169[7]), .SP(LOGIC_CLOCK_enable_148), 
            .CK(LOGIC_CLOCK), .Q(\writeData[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam writeData_i0_i7.GSR = "DISABLED";
    CCU2D add_7189_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n13156), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n13142), 
          .CIN(n10069), .COUT(n10070));
    defparam add_7189_13.INIT0 = 16'h00ae;
    defparam add_7189_13.INIT1 = 16'h00ae;
    defparam add_7189_13.INJECT1_0 = "NO";
    defparam add_7189_13.INJECT1_1 = "NO";
    LUT4 PIC_addr_31__I_0_i17_3_lut_rep_254_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[16]_adj_9 ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[16] ), 
         .Z(n12280)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam PIC_addr_31__I_0_i17_3_lut_rep_254_4_lut_4_lut.init = 16'h3808;
    LUT4 i8596_2_lut_rep_196_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[18] ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(n1921), 
         .Z(n12222)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i8596_2_lut_rep_196_3_lut_4_lut_4_lut.init = 16'hfff4;
    LUT4 BUS_VALID_N_477_I_0_2_lut_rep_203_3_lut_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[18] ), 
         .B(\BUS_currGrantID[1] ), .C(\BUS_currGrantID[0] ), .D(n2025), 
         .Z(LOGIC_CLOCK_enable_26)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam BUS_VALID_N_477_I_0_2_lut_rep_203_3_lut_4_lut_4_lut.init = 16'h000b;
    CCU2D add_7189_11 (.A0(\BUS_ADDR_INTERNAL[9] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13144), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n13143), 
          .CIN(n10068), .COUT(n10069));
    defparam add_7189_11.INIT0 = 16'h00dc;
    defparam add_7189_11.INIT1 = 16'hff51;
    defparam add_7189_11.INJECT1_0 = "NO";
    defparam add_7189_11.INJECT1_1 = "NO";
    FD1S3DX state_i1 (.D(state_7__N_1050[1]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_997), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i1.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_253_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[2] ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[2]_adj_15 ), .Z(n12279)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_253_4_lut_4_lut.init = 16'h3808;
    LUT4 i1_3_lut_rep_252_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[4] ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[4]_adj_16 ), .Z(n12278)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_252_4_lut_4_lut.init = 16'h3808;
    CCU2D add_7189_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[7]_adj_12 ), .D0(n13147), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), .D1(n13154), 
          .CIN(n10067), .COUT(n10068));
    defparam add_7189_9.INIT0 = 16'h00ae;
    defparam add_7189_9.INIT1 = 16'hff51;
    defparam add_7189_9.INJECT1_0 = "NO";
    defparam add_7189_9.INJECT1_1 = "NO";
    FD1P3DX state_i2 (.D(n13160), .SP(LOGIC_CLOCK_enable_149), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_997), .Q(state_c[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i2.GSR = "DISABLED";
    FD1P3DX state_i3 (.D(n13160), .SP(LOGIC_CLOCK_enable_150), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_997), .Q(state_c[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i3.GSR = "DISABLED";
    FD1S3DX state_i4 (.D(state_7__N_1050[4]), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_997), 
            .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i4.GSR = "DISABLED";
    FD1P3DX state_i5 (.D(n13160), .SP(LOGIC_CLOCK_enable_151), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_997), .Q(state_c[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i5.GSR = "DISABLED";
    FD1P3DX state_i6 (.D(n13160), .SP(LOGIC_CLOCK_enable_152), .CK(LOGIC_CLOCK), 
            .CD(BUS_DIRECTION_INTERNAL_N_997), .Q(state_c[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i6.GSR = "DISABLED";
    FD1S3DX state_i7 (.D(\state_7__N_1050[7] ), .CK(LOGIC_CLOCK), .CD(BUS_DIRECTION_INTERNAL_N_997), 
            .Q(\state[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam state_i7.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i1 (.D(data[9]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i1.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i2 (.D(data[10]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i2.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i3 (.D(data[11]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i3.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i4 (.D(data[12]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i4.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i5 (.D(data[13]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i5.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i6 (.D(data[14]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i6.GSR = "DISABLED";
    FD1P3AX rModDataTrans_i0_i7 (.D(data[15]), .SP(LOGIC_CLOCK_enable_159), 
            .CK(LOGIC_CLOCK), .Q(rModDataTrans[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=21, LSE_RCOL=36, LSE_LLINE=211, LSE_RLINE=211 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam rModDataTrans_i0_i7.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_247_4_lut_4_lut (.A(\BUS_ADDR_INTERNAL[8]_adj_1 ), .B(\BUS_currGrantID[1] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[8] ), .Z(n12273)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_3_lut_rep_247_4_lut_4_lut.init = 16'h3808;
    CCU2D add_7189_7 (.A0(\BUS_ADDR_INTERNAL[5]_adj_10 ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13145), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[6]_adj_11 ), 
          .D1(n13146), .CIN(n10066), .COUT(n10067));
    defparam add_7189_7.INIT0 = 16'h00dc;
    defparam add_7189_7.INIT1 = 16'h00ae;
    defparam add_7189_7.INJECT1_0 = "NO";
    defparam add_7189_7.INJECT1_1 = "NO";
    CCU2D add_7189_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[3]_adj_13 ), .D0(n13148), .A1(\BUS_ADDR_INTERNAL[4]_adj_16 ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13153), 
          .CIN(n10065), .COUT(n10066));
    defparam add_7189_5.INIT0 = 16'h00ae;
    defparam add_7189_5.INIT1 = 16'h00dc;
    defparam add_7189_5.INJECT1_0 = "NO";
    defparam add_7189_5.INJECT1_1 = "NO";
    CCU2D add_7189_3 (.A0(\BUS_ADDR_INTERNAL[1]_adj_14 ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13149), .A1(\BUS_ADDR_INTERNAL[2]_adj_15 ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13152), 
          .CIN(n10064), .COUT(n10065));
    defparam add_7189_3.INIT0 = 16'h00dc;
    defparam add_7189_3.INIT1 = 16'h00dc;
    defparam add_7189_3.INJECT1_0 = "NO";
    defparam add_7189_3.INJECT1_1 = "NO";
    CCU2D add_7189_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[0]_adj_17 ), 
          .D1(n12299), .COUT(n10064));
    defparam add_7189_1.INIT0 = 16'hF000;
    defparam add_7189_1.INIT1 = 16'h00ae;
    defparam add_7189_1.INJECT1_0 = "NO";
    defparam add_7189_1.INJECT1_1 = "NO";
    LUT4 mux_481_i2_4_lut (.A(rModDataWrite[9]), .B(PIC_DATA_IN_out_1), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i2_4_lut.init = 16'h0aca;
    LUT4 mux_481_i3_4_lut (.A(rModDataWrite[10]), .B(PIC_DATA_IN_out_2), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i3_4_lut.init = 16'h0aca;
    LUT4 mux_481_i4_4_lut (.A(rModDataWrite[11]), .B(PIC_DATA_IN_out_3), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i4_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_4_lut (.A(state[4]), .B(n12267), .C(\BUS_req[2] ), .D(n26), 
         .Z(n28)) /* synthesis lut_function=(A (D)+!A (B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut_4_lut.init = 16'hff45;
    LUT4 mux_481_i5_4_lut (.A(rModDataWrite[12]), .B(PIC_DATA_IN_out_4), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i5_4_lut.init = 16'h0aca;
    LUT4 mux_481_i6_4_lut (.A(rModDataWrite[13]), .B(PIC_DATA_IN_out_5), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i6_4_lut.init = 16'h0aca;
    LUT4 BUS_VALID_I_0_305_2_lut_rep_197 (.A(BUS_VALID_N_1118), .B(n2198), 
         .Z(n12223)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam BUS_VALID_I_0_305_2_lut_rep_197.init = 16'h2222;
    LUT4 i8686_2_lut_3_lut_4_lut (.A(BUS_VALID_N_1118), .B(n2198), .C(n13141), 
         .D(n19), .Z(LOGIC_CLOCK_enable_116)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam i8686_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i8707_3_lut_4_lut (.A(BUS_VALID_N_1118), .B(n2198), .C(n11485), 
         .D(n12219), .Z(LOGIC_CLOCK_enable_48)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(63[28:88])
    defparam i8707_3_lut_4_lut.init = 16'hd000;
    LUT4 mux_481_i7_4_lut (.A(rModDataWrite[14]), .B(PIC_DATA_IN_out_6), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i7_4_lut.init = 16'h0aca;
    LUT4 mux_481_i8_4_lut (.A(rModDataWrite[15]), .B(PIC_DATA_IN_out_7), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i8_4_lut.init = 16'h0aca;
    LUT4 i8587_4_lut (.A(n7167), .B(state_c[0]), .C(n38), .D(n12266), 
         .Z(state_7__N_1050[1])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i8587_4_lut.init = 16'h5f5d;
    LUT4 i1_3_lut_4_lut (.A(state[4]), .B(n12267), .C(n4_adj_1271), .D(state_c[0]), 
         .Z(n10891)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut (.A(n7167), .B(n12213), .C(state_c[2]), .D(n12293), 
         .Z(LOGIC_CLOCK_enable_149)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut.init = 16'h55d5;
    LUT4 readData_15__I_0_i3_4_lut (.A(n19), .B(writeData[2]), .C(n12314), 
         .D(transferMode[2]), .Z(\BUS_DATA_INTERNAL[2] )) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(68[23:106])
    defparam readData_15__I_0_i3_4_lut.init = 16'h5c0c;
    LUT4 i1_4_lut_adj_131 (.A(n7167), .B(n11014), .C(state_c[3]), .D(n12213), 
         .Z(LOGIC_CLOCK_enable_150)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut_adj_131.init = 16'h7555;
    LUT4 i1_2_lut_rep_210_3_lut_4_lut (.A(state[4]), .B(n12267), .C(PIC_WE_IN_c), 
         .D(state_c[0]), .Z(n12236)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_2_lut_rep_210_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_4_lut_adj_132 (.A(state[4]), .B(n23), .C(state[1]), .D(n12266), 
         .Z(state_7__N_1050[4])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut_adj_132.init = 16'heece;
    LUT4 i1_4_lut_adj_133 (.A(n7167), .B(state_c[5]), .C(n6), .D(state_c[3]), 
         .Z(LOGIC_CLOCK_enable_151)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut_adj_133.init = 16'h55d5;
    LUT4 i1_4_lut_adj_134 (.A(n7167), .B(n12213), .C(state_c[6]), .D(n11006), 
         .Z(LOGIC_CLOCK_enable_152)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut_adj_134.init = 16'h55d5;
    LUT4 i4815_2_lut (.A(PIC_DATA_IN_out_9), .B(PIC_WE_IN_c), .Z(data[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4815_2_lut.init = 16'h2222;
    LUT4 i4817_2_lut (.A(PIC_DATA_IN_out_11), .B(PIC_WE_IN_c), .Z(data[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4817_2_lut.init = 16'h2222;
    LUT4 i4818_2_lut (.A(PIC_DATA_IN_out_12), .B(PIC_WE_IN_c), .Z(data[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4818_2_lut.init = 16'h2222;
    LUT4 i4819_2_lut (.A(PIC_DATA_IN_out_13), .B(PIC_WE_IN_c), .Z(data[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4819_2_lut.init = 16'h2222;
    LUT4 i4820_2_lut (.A(PIC_DATA_IN_out_14), .B(PIC_WE_IN_c), .Z(data[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4820_2_lut.init = 16'h2222;
    LUT4 i4821_2_lut (.A(PIC_DATA_IN_out_15), .B(PIC_WE_IN_c), .Z(data[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4821_2_lut.init = 16'h2222;
    LUT4 i1_2_lut (.A(\BUS_req[2] ), .B(\BUS_currGrantID_3__N_72[0] ), .Z(\BUS_currGrantID_3__N_72[1] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut.init = 16'h2222;
    PFUMX i9055 (.BLUT(n12350), .ALUT(n12351), .C0(\BUS_currGrantID[1] ), 
          .Z(n12352));
    LUT4 i6_4_lut (.A(n11), .B(n12266), .C(n71), .D(\BUS_currGrantID[0] ), 
         .Z(LOGIC_CLOCK_enable_141)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i6_4_lut.init = 16'h0020;
    LUT4 i2_3_lut (.A(state_c[0]), .B(state[4]), .C(state[1]), .Z(n71)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i2_3_lut.init = 16'h0808;
    LUT4 PIC_OE_IN_I_0_2_lut_rep_319 (.A(PIC_OE_c), .B(PIC_WE_IN_c), .Z(n12345)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam PIC_OE_IN_I_0_2_lut_rep_319.init = 16'h8888;
    LUT4 BUS_DIRECTION_INTERNAL_I_105_2_lut_3_lut (.A(PIC_OE_c), .B(PIC_WE_IN_c), 
         .C(BUS_DIRECTION_INTERNAL_N_1000), .Z(BUS_DIRECTION_INTERNAL_N_997)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam BUS_DIRECTION_INTERNAL_I_105_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i8639_2_lut_3_lut (.A(PIC_OE_c), .B(PIC_WE_IN_c), .C(BUS_DIRECTION_INTERNAL_N_1000), 
         .Z(n11418)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[7:46])
    defparam i8639_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_320 (.A(state_c[6]), .B(\state[7] ), .Z(n12346)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_320.init = 16'heeee;
    LUT4 i8127_2_lut_3_lut_4_lut (.A(state_c[6]), .B(\state[7] ), .C(state_c[5]), 
         .D(state_c[2]), .Z(n11014)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i8127_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_286_3_lut (.A(state_c[6]), .B(\state[7] ), .C(state_c[2]), 
         .Z(n12312)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_286_3_lut.init = 16'hfefe;
    LUT4 i8694_2_lut_rep_297_3_lut (.A(state_c[6]), .B(\state[7] ), .C(state_c[5]), 
         .Z(n12323)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i8694_2_lut_rep_297_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_rep_267_3_lut_4_lut (.A(state_c[6]), .B(\state[7] ), .C(state_c[3]), 
         .D(state_c[5]), .Z(n12293)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_2_lut_rep_267_3_lut_4_lut.init = 16'hfffe;
    LUT4 i8637_4_lut (.A(n28), .B(n12293), .C(state[1]), .D(state_c[2]), 
         .Z(BUS_REQ_N_1209)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i8637_4_lut.init = 16'hfffd;
    LUT4 i8181_3_lut_4_lut_else_3_lut (.A(n12292), .B(\BUS_ADDR_INTERNAL[13] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_ADDR_INTERNAL[0]_adj_17 ), .Z(n12350)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C))) */ ;
    defparam i8181_3_lut_4_lut_else_3_lut.init = 16'he0c0;
    LUT4 i1_4_lut_adj_135 (.A(state_c[0]), .B(\BUS_req[2] ), .C(n12246), 
         .D(n12214), .Z(n26)) /* synthesis lut_function=(A ((C (D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i1_4_lut_adj_135.init = 16'ha222;
    LUT4 i1_2_lut_rep_321 (.A(state_c[2]), .B(state_c[3]), .Z(n12347)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_321.init = 16'heeee;
    LUT4 i8119_3_lut_4_lut (.A(state_c[2]), .B(state_c[3]), .C(state_c[5]), 
         .D(\state[7] ), .Z(n11006)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8119_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_298_3_lut (.A(state_c[2]), .B(state_c[3]), .C(state[1]), 
         .Z(n12324)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_298_3_lut.init = 16'hfefe;
    LUT4 i8640_4_lut (.A(n12246), .B(n11418), .C(n10258), .D(n15), .Z(LOGIC_CLOCK_enable_148)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;
    defparam i8640_4_lut.init = 16'h40c0;
    LUT4 mux_481_i1_4_lut (.A(rModDataWrite[8]), .B(PIC_DATA_IN_out_0), 
         .C(n15), .D(n12236), .Z(writeData_15__N_1169[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_481_i1_4_lut.init = 16'h0aca;
    LUT4 i4958_2_lut_rep_219_3_lut_4_lut (.A(state_c[3]), .B(n12323), .C(state[1]), 
         .D(state_c[2]), .Z(n12245)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(101[3] 156[10])
    defparam i4958_2_lut_rep_219_3_lut_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_adj_136 (.A(state[4]), .B(n7167), .Z(n15)) /* synthesis lut_function=((B)+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(125[10:23])
    defparam i1_2_lut_adj_136.init = 16'hdddd;
    LUT4 i1_2_lut_rep_213_3_lut_4_lut_4_lut (.A(n12323), .B(state[4]), .C(state_c[0]), 
         .D(n12324), .Z(n12239)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_2_lut_rep_213_3_lut_4_lut_4_lut.init = 16'hffdf;
    LUT4 i3_4_lut (.A(n12347), .B(n12323), .C(state_c[0]), .D(state[1]), 
         .Z(n7167)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i3_4_lut.init = 16'hfbff;
    LUT4 i8581_4_lut (.A(n7167), .B(n12245), .C(state_c[0]), .D(n12212), 
         .Z(state_7__N_1050[0])) /* synthesis lut_function=((B (C)+!B !(C (D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i8581_4_lut.init = 16'hd7f7;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\BUS_ADDR_INTERNAL[0] ), .B(n12348), .C(n12292), 
         .D(n13139), .Z(n6_adj_18)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    LUT4 i4814_2_lut (.A(PIC_DATA_IN_out_8), .B(PIC_WE_IN_c), .Z(data[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4814_2_lut.init = 16'h2222;
    LUT4 i4810_2_lut (.A(PIC_DATA_IN_out_4), .B(PIC_WE_IN_c), .Z(data[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4810_2_lut.init = 16'h2222;
    CCU2D lastAddress_18__I_0_19 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n9697), .S0(BUS_DIRECTION_INTERNAL_N_1000));
    defparam lastAddress_18__I_0_19.INIT0 = 16'hFFFF;
    defparam lastAddress_18__I_0_19.INIT1 = 16'h0000;
    defparam lastAddress_18__I_0_19.INJECT1_0 = "NO";
    defparam lastAddress_18__I_0_19.INJECT1_1 = "NO";
    LUT4 readData_15__I_0_i2_4_lut (.A(n19), .B(writeData[1]), .C(n12314), 
         .D(transferMode[1]), .Z(\BUS_DATA_INTERNAL[1] )) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(68[23:106])
    defparam readData_15__I_0_i2_4_lut.init = 16'h5c0c;
    LUT4 i1_4_lut_adj_137 (.A(transferMode[0]), .B(transferMode[1]), .C(transferMode[2]), 
         .D(n10324), .Z(n23_adj_1273)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_137.init = 16'h0002;
    LUT4 i8_4_lut (.A(data[10]), .B(n16), .C(PIC_DATA_IN_out_12), .D(PIC_DATA_IN_out_11), 
         .Z(n10324)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i7_4_lut (.A(PIC_DATA_IN_out_13), .B(PIC_DATA_IN_out_15), .C(PIC_DATA_IN_out_9), 
         .D(n10), .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_138 (.A(PIC_DATA_IN_out_8), .B(PIC_DATA_IN_out_14), 
         .Z(n10)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i1_2_lut_adj_138.init = 16'h8888;
    LUT4 i2_2_lut (.A(PIC_DATA_IN_out_10), .B(PIC_WE_IN_c), .Z(data[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i2_2_lut.init = 16'h2222;
    LUT4 i8181_3_lut_4_lut_then_3_lut (.A(n12292), .B(\BUS_currGrantID[0] ), 
         .C(\BUS_ADDR_INTERNAL[0] ), .Z(n12351)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i8181_3_lut_4_lut_then_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_139 (.A(n10895), .B(n12273), .C(n69), 
         .D(n5045), .Z(n1184)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_2_lut_3_lut_4_lut_adj_139.init = 16'hfffd;
    LUT4 i6492_4_lut (.A(\BUS_currGrantID[1] ), .B(\BUS_currGrantID_3__N_72[0] ), 
         .C(\BUS_currGrantID[0] ), .D(\BUS_req[2] ), .Z(BUS_currGrantID_3__N_54)) /* synthesis lut_function=(A (C+!(D))+!A !(B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(56[8:23])
    defparam i6492_4_lut.init = 16'hb0ba;
    LUT4 i2737_3_lut_4_lut (.A(PIC_WE_IN_c), .B(n12239), .C(n15), .D(LOGIC_CLOCK_enable_148), 
         .Z(n5334)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i2737_3_lut_4_lut.init = 16'hef00;
    LUT4 i4_3_lut_4_lut (.A(BUS_DIRECTION_INTERNAL_N_1000), .B(n12345), 
         .C(\BUS_currGrantID[1] ), .D(BUS_DONE), .Z(n11)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i4_3_lut_4_lut.init = 16'h2000;
    LUT4 n23_bdd_3_lut (.A(n23_adj_1273), .B(transferMode[3]), .C(PIC_WE_IN_c), 
         .Z(n11759)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n23_bdd_3_lut.init = 16'h0202;
    LUT4 i1_4_lut_adj_140 (.A(state[4]), .B(PIC_WE_IN_c), .C(n8), .D(state_c[3]), 
         .Z(n14)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_4_lut_adj_140.init = 16'haaba;
    LUT4 i3328_4_lut (.A(transferMode[0]), .B(writeData[0]), .C(n12314), 
         .D(n19), .Z(\BUS_DATA_INTERNAL[0] )) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(39[8:25])
    defparam i3328_4_lut.init = 16'h0cac;
    LUT4 i3_4_lut_adj_141 (.A(n5045), .B(n12250), .C(n10895), .D(n69), 
         .Z(n19)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i3_4_lut_adj_141.init = 16'hffbf;
    LUT4 i2_2_lut_3_lut_4_lut (.A(n12246), .B(state_c[0]), .C(n12345), 
         .D(BUS_DIRECTION_INTERNAL_N_1000), .Z(LOGIC_CLOCK_enable_159)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i4863_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[9]), .D(n12217), .Z(\PIC_data[9] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4863_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4865_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[11]), .D(n12217), .Z(\PIC_data[11] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4865_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4864_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[10]), .D(n12217), .Z(\PIC_data[10] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4864_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i104_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[15]), .D(n12217), .Z(n100)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i104_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4866_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[12]), .D(n12217), .Z(\PIC_data[12] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4866_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4862_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[8]), .D(n12217), .Z(\PIC_data[8] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4862_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4867_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[13]), .D(n12217), .Z(\PIC_data[13] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4867_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i4868_2_lut_3_lut_4_lut (.A(n12348), .B(BUS_DIRECTION_INTERNAL), 
         .C(writeData[14]), .D(n12217), .Z(\PIC_data[14] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4868_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 lastAddress_i1_i5_3_lut_4_lut (.A(n12344), .B(n12278), .C(SRAM_WE_N_704), 
         .D(\lastAddress[4] ), .Z(n60)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam lastAddress_i1_i5_3_lut_4_lut.init = 16'hfd0d;
    LUT4 i1_4_lut_adj_142 (.A(n12214), .B(state[1]), .C(n12266), .D(state_c[0]), 
         .Z(LOGIC_CLOCK_enable_46)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/sram.vhd(34[8:13])
    defparam i1_4_lut_adj_142.init = 16'ha8a0;
    LUT4 i3_4_lut_adj_143 (.A(state_c[0]), .B(n10904), .C(n12323), .D(n11418), 
         .Z(LOGIC_CLOCK_enable_47)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_143.init = 16'h8000;
    LUT4 i1_4_lut_adj_144 (.A(PIC_WE_IN_c), .B(state[4]), .C(n12242), 
         .D(n12267), .Z(n4_adj_1271)) /* synthesis lut_function=(A ((D)+!B)+!A (B (C (D))+!B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    defparam i1_4_lut_adj_144.init = 16'hfa32;
    CCU2D lastAddress_18__I_0_19_7181 (.A0(PIC_ADDR_IN_c_3), .B0(lastAddress[3]), 
          .C0(PIC_ADDR_IN_c_2), .D0(lastAddress[2]), .A1(PIC_ADDR_IN_c_1), 
          .B1(lastAddress[1]), .C1(PIC_ADDR_IN_c_0), .D1(lastAddress[0]), 
          .CIN(n9696), .COUT(n9697));
    defparam lastAddress_18__I_0_19_7181.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_19_7181.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_19_7181.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_19_7181.INJECT1_1 = "YES";
    LUT4 lastAddress_i1_i8_3_lut_3_lut_4_lut (.A(n12344), .B(n12288), .C(\lastAddress[7] ), 
         .D(SRAM_WE_N_704), .Z(n57)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C+!(D))) */ ;
    defparam lastAddress_i1_i8_3_lut_3_lut_4_lut.init = 16'hf0dd;
    LUT4 lastAddress_i1_i4_3_lut_4_lut (.A(n12344), .B(n12287), .C(SRAM_WE_N_704), 
         .D(\lastAddress[3] ), .Z(n61)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam lastAddress_i1_i4_3_lut_4_lut.init = 16'hfd0d;
    LUT4 i2_3_lut_4_lut_adj_145 (.A(state_c[5]), .B(n12346), .C(n12347), 
         .D(state[1]), .Z(n4)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i2_3_lut_4_lut_adj_145.init = 16'h0100;
    LUT4 i1_2_lut_rep_240_3_lut_4_lut (.A(state_c[5]), .B(n12346), .C(state_c[2]), 
         .D(state_c[3]), .Z(n12266)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_2_lut_rep_240_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_220_3_lut_3_lut_4_lut (.A(state_c[5]), .B(n12346), 
         .C(n12324), .D(state[4]), .Z(n12246)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_2_lut_rep_220_3_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_241_2_lut_3_lut_4_lut (.A(state[1]), .B(n12347), .C(n12346), 
         .D(state_c[5]), .Z(n12267)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_241_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_146 (.A(state_c[2]), .B(n12293), .C(n11760), 
         .D(state[1]), .Z(n38)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(108[4] 154[11])
    defparam i1_3_lut_4_lut_adj_146.init = 16'h00fe;
    LUT4 lastAddress_i1_i18_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(SRAM_WE_N_704), 
         .C(\lastAddress[17] ), .D(n13158), .Z(n47)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A ((C)+!B)) */ ;
    defparam lastAddress_i1_i18_3_lut_3_lut_4_lut_4_lut.init = 16'hd1f3;
    LUT4 i1_2_lut_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n12344), .B(n13158), 
         .C(n13140), .D(n12304), .Z(lastAddress_31__N_833)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_2_lut_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h8880;
    LUT4 i1_2_lut_2_lut_3_lut_3_lut_4_lut_4_lut_adj_147 (.A(n12344), .B(n13158), 
         .C(n13140), .D(n12304), .Z(lastAddress_31__N_773)) /* synthesis lut_function=(!(A (B+!(C+(D))))) */ ;
    defparam i1_2_lut_2_lut_3_lut_3_lut_4_lut_4_lut_adj_147.init = 16'h7775;
    LUT4 i7296_4_lut_4_lut_4_lut_4_lut (.A(n12344), .B(n13158), .C(n9924), 
         .D(n12304), .Z(BUS_DONE_OUT_N_626)) /* synthesis lut_function=((B (C (D))+!B (D))+!A) */ ;
    defparam i7296_4_lut_4_lut_4_lut_4_lut.init = 16'hf755;
    LUT4 readData_15__I_0_i4_4_lut (.A(transferMode[3]), .B(writeData[3]), 
         .C(n12314), .D(n19), .Z(\BUS_DATA_INTERNAL[3] )) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(68[23:106])
    defparam readData_15__I_0_i4_4_lut.init = 16'h0cac;
    CCU2D lastAddress_18__I_0_17 (.A0(PIC_ADDR_IN_c_7), .B0(lastAddress[7]), 
          .C0(PIC_ADDR_IN_c_6), .D0(lastAddress[6]), .A1(PIC_ADDR_IN_c_5), 
          .B1(lastAddress[5]), .C1(PIC_ADDR_IN_c_4), .D1(lastAddress[4]), 
          .CIN(n9695), .COUT(n9696));
    defparam lastAddress_18__I_0_17.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_17.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_17.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_17.INJECT1_1 = "YES";
    LUT4 i1_2_lut_rep_216 (.A(n23_adj_1273), .B(transferMode[3]), .Z(n12242)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    defparam i1_2_lut_rep_216.init = 16'h2222;
    LUT4 i3_3_lut_4_lut (.A(n23_adj_1273), .B(transferMode[3]), .C(state[1]), 
         .D(n11014), .Z(n8)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(24[3:12])
    defparam i3_3_lut_4_lut.init = 16'h0002;
    CCU2D lastAddress_18__I_0_15 (.A0(PIC_ADDR_IN_c_11), .B0(lastAddress[11]), 
          .C0(PIC_ADDR_IN_c_10), .D0(lastAddress[10]), .A1(PIC_ADDR_IN_c_9), 
          .B1(lastAddress[9]), .C1(PIC_ADDR_IN_c_8), .D1(lastAddress[8]), 
          .CIN(n9694), .COUT(n9695));
    defparam lastAddress_18__I_0_15.INIT0 = 16'h9009;
    defparam lastAddress_18__I_0_15.INIT1 = 16'h9009;
    defparam lastAddress_18__I_0_15.INJECT1_0 = "YES";
    defparam lastAddress_18__I_0_15.INJECT1_1 = "YES";
    CCU2D add_313_9 (.A0(rModDataTrans[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10019), .S0(rModDataWrite_15__N_1120[7]), .S1(rModDataWrite_15__N_1120[8]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_313_9.INIT0 = 16'hf555;
    defparam add_313_9.INIT1 = 16'h0000;
    defparam add_313_9.INJECT1_0 = "NO";
    defparam add_313_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_207_4_lut (.A(n13154), .B(\BUS_ADDR_INTERNAL[8] ), 
         .C(n12332), .D(n10895), .Z(n12233)) /* synthesis lut_function=(A+!(B (C (D))+!B (D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(67[18:73])
    defparam i1_2_lut_rep_207_4_lut.init = 16'haeff;
    CCU2D add_313_7 (.A0(rModDataTrans[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(rModDataTrans[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10018), .COUT(n10019), .S0(rModDataWrite_15__N_1120[5]), 
          .S1(rModDataWrite_15__N_1120[6]));   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(94[63:82])
    defparam add_313_7.INIT0 = 16'hf555;
    defparam add_313_7.INIT1 = 16'hf555;
    defparam add_313_7.INJECT1_0 = "NO";
    defparam add_313_7.INJECT1_1 = "NO";
    LUT4 i4623_2_lut (.A(PIC_DATA_IN_out_0), .B(PIC_WE_IN_c), .Z(data[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4623_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_4_lut (.A(\BUS_ADDR_INTERNAL[4]_adj_16 ), .B(n13153), 
         .C(n12332), .D(n12287), .Z(n10976)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam i1_2_lut_4_lut.init = 16'hffce;
    LUT4 i4808_2_lut (.A(PIC_DATA_IN_out_2), .B(PIC_WE_IN_c), .Z(data[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4808_2_lut.init = 16'h2222;
    LUT4 i8125_2_lut_4_lut (.A(\BUS_ADDR_INTERNAL[4]_adj_16 ), .B(n13153), 
         .C(n12332), .D(n12279), .Z(n11012)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(105[14:81])
    defparam i8125_2_lut_4_lut.init = 16'hffce;
    LUT4 i4807_2_lut (.A(PIC_DATA_IN_out_1), .B(PIC_WE_IN_c), .Z(data[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/pic.vhd(98[10:55])
    defparam i4807_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module MatrixDriver
//

module MatrixDriver (PIXEL_CLOCK, \BUS_currGrantID[0] , \BUS_currGrantID[1] , 
            GND_net, BUS_VALID_N_113, Matrix_LINE_SEL_Out_c_0, \BUS_ADDR_INTERNAL[18] , 
            n12309, Matrix_CTRL_Out_c_1, PIXEL_CLOCK_N_302, \BUS_ADDR_INTERNAL[16] , 
            n13151, n13158, n12344, currPWMCount, LOGIC_CLOCK, \BUS_ADDR_INTERNAL[14] , 
            n13157, \BUS_ADDR_INTERNAL[15] , n13150, WRITE_DONE, LOGIC_CLOCK_N_116, 
            PWMArray_0__12__N_110, n13160, \PWMArray[0][12] , \BUS_data[3] , 
            \currPWMCountMax[0] , \BUS_ADDR_INTERNAL[12] , n13142, \BUS_ADDR_INTERNAL[13] , 
            n13155, \BUS_ADDR_INTERNAL[10] , n13143, \BUS_ADDR_INTERNAL[11] , 
            n13156, \PWMArray[0][11] , \BUS_data[2] , \BUS_ADDR_INTERNAL[8] , 
            n13154, \BUS_ADDR_INTERNAL[9] , n13144, \BUS_ADDR_INTERNAL[7] , 
            n13147, MATRIX_CURRROW, \PWMArray[0][9] , \BUS_data[0] , 
            \PWMArray[0][10] , \BUS_data[1] , \currPWMCountMax[2] , \currPWMCountMax[5] , 
            \currPWMCountMax[1] , \currPWMCountMax[4] , \currPWMCountMax[3] , 
            \currPWMCountMax[6] , Matrix_LINE_SEL_Out_c_1, n1886, \currPWMCountMax[12] , 
            Matrix_CTRL_Out_c_2, \currPWMCountMax[11] , \currPWMCountMax[10] , 
            \currPWMCountMax[9] , \currPWMCountMax[8] , \currPWMCountMax[7] , 
            \BUS_ADDR_INTERNAL[5] , n13145, \BUS_ADDR_INTERNAL[6] , n13146, 
            \BUS_ADDR_INTERNAL[3] , n13148, \BUS_ADDR_INTERNAL[4] , n13153, 
            \BUS_ADDR_INTERNAL[1] , n13149, \BUS_ADDR_INTERNAL[2] , n13152, 
            \BUS_ADDR_INTERNAL[0] , n12299, currReadRow, n12231, Matrix_DATA_Out_c_11, 
            Matrix_DATA_Out_c_10, Matrix_DATA_Out_c_9, Matrix_DATA_Out_c_8, 
            Matrix_DATA_Out_c_7, Matrix_DATA_Out_c_6, Matrix_DATA_Out_c_5, 
            Matrix_DATA_Out_c_4, Matrix_DATA_Out_c_3, Matrix_DATA_Out_c_2, 
            Matrix_DATA_Out_c_1, Matrix_DATA_Out_c_0, Matrix_LINE_SEL_Out_c_2, 
            Matrix_CTRL_Out_c_0, n12311, \lastReadRow[4] , n10349, n12221, 
            n13141, n87, \lastReadRow[3] , n12342, n10350, n12284, 
            \VRAM_ADDR[6] , \VRAM_ADDR[5] , \VRAM_ADDR[4] , \VRAM_ADDR[3] , 
            \VRAM_ADDR[2] , \VRAM_ADDR[1] , \VRAM_ADDR[0] , n3028, n3027, 
            VCC_net, VRAM_WC, n3035, n3034, n3033, n3032, n3037, 
            n3036, n3030, n3029, n3031, VRAM_DATA);
    input PIXEL_CLOCK;
    input \BUS_currGrantID[0] ;
    input \BUS_currGrantID[1] ;
    input GND_net;
    output BUS_VALID_N_113;
    output Matrix_LINE_SEL_Out_c_0;
    input \BUS_ADDR_INTERNAL[18] ;
    input n12309;
    output Matrix_CTRL_Out_c_1;
    input PIXEL_CLOCK_N_302;
    input \BUS_ADDR_INTERNAL[16] ;
    input n13151;
    input n13158;
    input n12344;
    output [15:0]currPWMCount;
    input LOGIC_CLOCK;
    input \BUS_ADDR_INTERNAL[14] ;
    input n13157;
    input \BUS_ADDR_INTERNAL[15] ;
    input n13150;
    output WRITE_DONE;
    input LOGIC_CLOCK_N_116;
    input PWMArray_0__12__N_110;
    input n13160;
    output \PWMArray[0][12] ;
    input \BUS_data[3] ;
    output \currPWMCountMax[0] ;
    input \BUS_ADDR_INTERNAL[12] ;
    input n13142;
    input \BUS_ADDR_INTERNAL[13] ;
    input n13155;
    input \BUS_ADDR_INTERNAL[10] ;
    input n13143;
    input \BUS_ADDR_INTERNAL[11] ;
    input n13156;
    output \PWMArray[0][11] ;
    input \BUS_data[2] ;
    input \BUS_ADDR_INTERNAL[8] ;
    input n13154;
    input \BUS_ADDR_INTERNAL[9] ;
    input n13144;
    input \BUS_ADDR_INTERNAL[7] ;
    input n13147;
    output [4:0]MATRIX_CURRROW;
    output \PWMArray[0][9] ;
    input \BUS_data[0] ;
    output \PWMArray[0][10] ;
    input \BUS_data[1] ;
    output \currPWMCountMax[2] ;
    output \currPWMCountMax[5] ;
    output \currPWMCountMax[1] ;
    output \currPWMCountMax[4] ;
    output \currPWMCountMax[3] ;
    output \currPWMCountMax[6] ;
    output Matrix_LINE_SEL_Out_c_1;
    output n1886;
    output \currPWMCountMax[12] ;
    output Matrix_CTRL_Out_c_2;
    output \currPWMCountMax[11] ;
    output \currPWMCountMax[10] ;
    output \currPWMCountMax[9] ;
    output \currPWMCountMax[8] ;
    output \currPWMCountMax[7] ;
    input \BUS_ADDR_INTERNAL[5] ;
    input n13145;
    input \BUS_ADDR_INTERNAL[6] ;
    input n13146;
    input \BUS_ADDR_INTERNAL[3] ;
    input n13148;
    input \BUS_ADDR_INTERNAL[4] ;
    input n13153;
    input \BUS_ADDR_INTERNAL[1] ;
    input n13149;
    input \BUS_ADDR_INTERNAL[2] ;
    input n13152;
    input \BUS_ADDR_INTERNAL[0] ;
    input n12299;
    output [4:0]currReadRow;
    input n12231;
    output Matrix_DATA_Out_c_11;
    output Matrix_DATA_Out_c_10;
    output Matrix_DATA_Out_c_9;
    output Matrix_DATA_Out_c_8;
    output Matrix_DATA_Out_c_7;
    output Matrix_DATA_Out_c_6;
    output Matrix_DATA_Out_c_5;
    output Matrix_DATA_Out_c_4;
    output Matrix_DATA_Out_c_3;
    output Matrix_DATA_Out_c_2;
    output Matrix_DATA_Out_c_1;
    output Matrix_DATA_Out_c_0;
    output Matrix_LINE_SEL_Out_c_2;
    output Matrix_CTRL_Out_c_0;
    output n12311;
    input \lastReadRow[4] ;
    output n10349;
    output n12221;
    input n13141;
    input n87;
    input \lastReadRow[3] ;
    output n12342;
    output n10350;
    output n12284;
    input \VRAM_ADDR[6] ;
    input \VRAM_ADDR[5] ;
    input \VRAM_ADDR[4] ;
    input \VRAM_ADDR[3] ;
    input \VRAM_ADDR[2] ;
    input \VRAM_ADDR[1] ;
    input \VRAM_ADDR[0] ;
    input [9:0]n3028;
    input [9:0]n3027;
    input VCC_net;
    input VRAM_WC;
    input [9:0]n3035;
    input [9:0]n3034;
    input [9:0]n3033;
    input [9:0]n3032;
    input [9:0]n3037;
    input [9:0]n3036;
    input [9:0]n3030;
    input [9:0]n3029;
    input [9:0]n3031;
    input [9:0]VRAM_DATA;
    
    wire PIXEL_CLOCK /* synthesis SET_AS_NETWORK=PIXEL_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(43[8:19])
    wire PIXEL_CLOCK_N_302 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(82[9:22])
    wire LOGIC_CLOCK /* synthesis SET_AS_NETWORK=LOGIC_CLOCK, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(44[8:19])
    wire LOGIC_CLOCK_N_116 /* synthesis is_clock=1, is_inv_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(73[9:17])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(90[8:15])
    
    wire n11286, n11287;
    wire [3:0]currBit;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(60[9:16])
    
    wire n11288, PIXEL_CLOCK_enable_13, PIXEL_CLOCK_enable_24, n12339, 
        n11293, n11294, n11295, n11300, n11301, n11302, n11307, 
        n11308, n11309, n10187, n11314, n11315, n11316, PIXEL_CLOCK_enable_2, 
        n12243, n11321, n11322, n11323, n10186, PIXEL_CLOCK_enable_3, 
        n2, n11240, n11241, n11244;
    wire [15:0]currPWMVal;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(85[9:19])
    
    wire PIXEL_CLOCK_N_302_enable_26;
    wire [15:0]currPWMVal_15__N_213;
    
    wire n10185, MATRIX_CLKEN_LAT, MATRIX_CLKEN, LOGIC_CLOCK_enable_64;
    wire [15:0]currPWMCount_15__N_149;
    
    wire n10184, LOGIC_CLOCK_N_116_enable_22, n7141, n12298, PIXEL_CLOCK_enable_4, 
        n12240, n11242, n11243, n11245, n10183, n10182, n11247, 
        n11248, n11251, n11249, n11250, n11252, n10181, n11254, 
        n11255, n11258, n11256, n11257, n11259;
    wire [7:0]VRAM_READ_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(79[9:23])
    
    wire VRAM_READ_ADDR_7__N_127, n11261, n11262, n11265, n28, n11263, 
        n11264, n11266, n11724, n12349;
    wire [15:0]currPWMCountMax_15__N_230;
    wire [7:0]currPixel;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(59[9:18])
    
    wire PIXEL_CLOCK_enable_25, n5345;
    wire [7:0]n37;
    
    wire n11268, n11269, n11272;
    wire [3:0]n21;
    
    wire n11270, n11271, n11273;
    wire [4:0]lastRow;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(62[9:16])
    
    wire PIXEL_CLOCK_enable_20, n11275, n11276, n11279;
    wire [4:0]n12;
    
    wire n5332, n3, n5322, n7, n3_adj_1219, n13137, n13138, n12333, 
        n7_adj_1220, n7_adj_1221, n9971;
    wire [15:0]currPWMCount_15__N_262;
    
    wire n9972, PIXEL_CLOCK_enable_15, n12254, n10116, n10115, n11303, 
        n11304, n10114, n10113, n10003, n10112, n10002, n10001, 
        n10111, n10000, n11277, n11278, n11280, n10110, n9999, 
        n10109, n22_adj_1222, n30, n10108, n10107, n11282, n11283, 
        n10106;
    wire [7:0]n47;
    
    wire n9998, n9997, n11284, n11285, n11289, n11290, n11291, 
        n11292, n9996, n11296, n11297, n11298, n11299;
    wire [9:0]\RED[1] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(68[9:12])
    
    wire n12260, n12249, n1095, n11246, n8;
    wire [9:0]\BLUE[3] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(70[9:13])
    
    wire n11253, n8_adj_1223;
    wire [9:0]\GREEN[3] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(69[9:14])
    
    wire n11260, n8_adj_1224;
    wire [9:0]\RED[3] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(68[9:12])
    
    wire n11267, n8_adj_1225;
    wire [9:0]\BLUE[2] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(70[9:13])
    
    wire n11274, n8_adj_1226, n10_adj_1227;
    wire [9:0]\GREEN[2] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(69[9:14])
    
    wire n11281, n8_adj_1228;
    wire [9:0]\RED[2] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(68[9:12])
    
    wire n8_adj_1229;
    wire [9:0]\BLUE[1] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(70[9:13])
    
    wire n8_adj_1230, n12306, n14;
    wire [9:0]\GREEN[1] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(69[9:14])
    
    wire n8_adj_1231, n8_adj_1232;
    wire [9:0]\BLUE[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(70[9:13])
    
    wire n8_adj_1233;
    wire [9:0]\GREEN[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(69[9:14])
    
    wire n8_adj_1234;
    wire [9:0]\RED[0] ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(68[9:12])
    
    wire n6, n11320, n11319, n11318, n12336, n12135, n11317, n11313, 
        n10037, n11312, n11311, n11310, n10036, n9970, n12334, 
        n12359, n12357, n10035, n10034, n12047, n9969, n12330, 
        n12275, MATRIX_ROWCLK_N_289, n11306, n11305;
    wire [7:0]VRAM_WRITE_ADDR;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(100[9:24])
    
    wire n12335, n12340, n7_adj_1235, n7_adj_1236, n12337, n26, 
        n25, n12285, n14_adj_1237, n12281, n11718, n7_adj_1238, 
        n6_adj_1239, n9975, n12241, n6_adj_1240, n11924, n9968, 
        n14_adj_1241, n9974, n9973;
    
    L6MUX21 i8396 (.D0(n11286), .D1(n11287), .SD(currBit[2]), .Z(n11288));
    FD1P3IX currBit_680__i0 (.D(n12339), .SP(PIXEL_CLOCK_enable_13), .CD(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(currBit[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_680__i0.GSR = "DISABLED";
    L6MUX21 i8403 (.D0(n11293), .D1(n11294), .SD(currBit[2]), .Z(n11295));
    L6MUX21 i8410 (.D0(n11300), .D1(n11301), .SD(currBit[2]), .Z(n11302));
    L6MUX21 i8417 (.D0(n11307), .D1(n11308), .SD(currBit[2]), .Z(n11309));
    CCU2D add_7183_15 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10187), .S1(BUS_VALID_N_113));
    defparam add_7183_15.INIT0 = 16'heeee;
    defparam add_7183_15.INIT1 = 16'h0000;
    defparam add_7183_15.INJECT1_0 = "NO";
    defparam add_7183_15.INJECT1_1 = "NO";
    L6MUX21 i8424 (.D0(n11314), .D1(n11315), .SD(currBit[2]), .Z(n11316));
    FD1P3AX MATRIX_ROWCLK_148 (.D(n12243), .SP(PIXEL_CLOCK_enable_2), .CK(PIXEL_CLOCK), 
            .Q(Matrix_LINE_SEL_Out_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam MATRIX_ROWCLK_148.GSR = "DISABLED";
    L6MUX21 i8431 (.D0(n11321), .D1(n11322), .SD(currBit[2]), .Z(n11323));
    CCU2D add_7183_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[18] ), .D0(n12309), .A1(\BUS_currGrantID[0] ), 
          .B1(\BUS_currGrantID[1] ), .C1(GND_net), .D1(GND_net), .CIN(n10186), 
          .COUT(n10187));
    defparam add_7183_13.INIT0 = 16'hff20;
    defparam add_7183_13.INIT1 = 16'heeee;
    defparam add_7183_13.INJECT1_0 = "NO";
    defparam add_7183_13.INJECT1_1 = "NO";
    FD1P3AX MATRIX_LAT_146 (.D(n2), .SP(PIXEL_CLOCK_enable_3), .CK(PIXEL_CLOCK), 
            .Q(Matrix_CTRL_Out_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam MATRIX_LAT_146.GSR = "DISABLED";
    PFUMX i8352 (.BLUT(n11240), .ALUT(n11241), .C0(currBit[1]), .Z(n11244));
    FD1P3AX currPWMVal_i0_i0 (.D(currPWMVal_15__N_213[0]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i0.GSR = "DISABLED";
    CCU2D add_7183_11 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[16] ), .D0(n13151), .A1(n13158), .B1(n12344), 
          .C1(GND_net), .D1(GND_net), .CIN(n10185), .COUT(n10186));
    defparam add_7183_11.INIT0 = 16'h00ae;
    defparam add_7183_11.INIT1 = 16'h8888;
    defparam add_7183_11.INJECT1_0 = "NO";
    defparam add_7183_11.INJECT1_1 = "NO";
    FD1S3AX MATRIX_CLKEN_LAT_155 (.D(MATRIX_CLKEN), .CK(PIXEL_CLOCK_N_302), 
            .Q(MATRIX_CLKEN_LAT)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam MATRIX_CLKEN_LAT_155.GSR = "DISABLED";
    FD1P3BX currPWMCount_i0 (.D(currPWMCount_15__N_149[0]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i0.GSR = "DISABLED";
    CCU2D add_7183_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[14] ), .D0(n13157), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[15] ), .D1(n13150), 
          .CIN(n10184), .COUT(n10185));
    defparam add_7183_9.INIT0 = 16'h00ae;
    defparam add_7183_9.INIT1 = 16'h00ae;
    defparam add_7183_9.INJECT1_0 = "NO";
    defparam add_7183_9.INJECT1_1 = "NO";
    FD1S3DX WRITE_DONE_158 (.D(n13160), .CK(LOGIC_CLOCK_N_116), .CD(PWMArray_0__12__N_110), 
            .Q(WRITE_DONE)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam WRITE_DONE_158.GSR = "DISABLED";
    FD1P3AY brightness_3__159 (.D(\BUS_data[3] ), .SP(LOGIC_CLOCK_N_116_enable_22), 
            .CK(LOGIC_CLOCK_N_116), .Q(\PWMArray[0][12] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam brightness_3__159.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i1 (.D(n12298), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n7141), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i1.GSR = "DISABLED";
    FD1P3IX MATRIX_CLKEN_145 (.D(n13160), .SP(PIXEL_CLOCK_enable_4), .CD(n12240), 
            .CK(PIXEL_CLOCK), .Q(MATRIX_CLKEN)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam MATRIX_CLKEN_145.GSR = "DISABLED";
    PFUMX i8353 (.BLUT(n11242), .ALUT(n11243), .C0(currBit[1]), .Z(n11245));
    CCU2D add_7183_7 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[12] ), .D0(n13142), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[13] ), .D1(n13155), 
          .CIN(n10183), .COUT(n10184));
    defparam add_7183_7.INIT0 = 16'h00ae;
    defparam add_7183_7.INIT1 = 16'h00ae;
    defparam add_7183_7.INJECT1_0 = "NO";
    defparam add_7183_7.INJECT1_1 = "NO";
    CCU2D add_7183_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[10] ), .D0(n13143), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[11] ), .D1(n13156), 
          .CIN(n10182), .COUT(n10183));
    defparam add_7183_5.INIT0 = 16'hff51;
    defparam add_7183_5.INIT1 = 16'h00ae;
    defparam add_7183_5.INJECT1_0 = "NO";
    defparam add_7183_5.INJECT1_1 = "NO";
    PFUMX i8359 (.BLUT(n11247), .ALUT(n11248), .C0(currBit[1]), .Z(n11251));
    FD1P3AY brightness_2__160 (.D(\BUS_data[2] ), .SP(LOGIC_CLOCK_N_116_enable_22), 
            .CK(LOGIC_CLOCK_N_116), .Q(\PWMArray[0][11] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam brightness_2__160.GSR = "DISABLED";
    PFUMX i8360 (.BLUT(n11249), .ALUT(n11250), .C0(currBit[1]), .Z(n11252));
    CCU2D add_7183_3 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[8] ), .D0(n13154), .A1(\BUS_ADDR_INTERNAL[9] ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13144), 
          .CIN(n10181), .COUT(n10182));
    defparam add_7183_3.INIT0 = 16'h00ae;
    defparam add_7183_3.INIT1 = 16'h00dc;
    defparam add_7183_3.INJECT1_0 = "NO";
    defparam add_7183_3.INJECT1_1 = "NO";
    CCU2D add_7183_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[7] ), 
          .D1(n13147), .COUT(n10181));
    defparam add_7183_1.INIT0 = 16'hF000;
    defparam add_7183_1.INIT1 = 16'h00ae;
    defparam add_7183_1.INJECT1_0 = "NO";
    defparam add_7183_1.INJECT1_1 = "NO";
    PFUMX i8366 (.BLUT(n11254), .ALUT(n11255), .C0(currBit[1]), .Z(n11258));
    PFUMX i8367 (.BLUT(n11256), .ALUT(n11257), .C0(currBit[1]), .Z(n11259));
    FD1P3AX VRAM_PAGEMAPPING_152 (.D(VRAM_READ_ADDR_7__N_127), .SP(PIXEL_CLOCK_enable_13), 
            .CK(PIXEL_CLOCK), .Q(VRAM_READ_ADDR[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam VRAM_PAGEMAPPING_152.GSR = "DISABLED";
    PFUMX i8373 (.BLUT(n11261), .ALUT(n11262), .C0(currBit[1]), .Z(n11265));
    LUT4 i12_4_lut (.A(currPWMCount[11]), .B(currPWMCount[9]), .C(currPWMCount[14]), 
         .D(currPWMCount[15]), .Z(n28)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut.init = 16'h8000;
    PFUMX i8374 (.BLUT(n11263), .ALUT(n11264), .C0(currBit[1]), .Z(n11266));
    PFUMX i8769 (.BLUT(n11724), .ALUT(n12349), .C0(currBit[3]), .Z(currPWMCountMax_15__N_230[9]));
    FD1P3IX currPixel_679__i6 (.D(n37[6]), .SP(PIXEL_CLOCK_enable_25), .CD(n5345), 
            .CK(PIXEL_CLOCK), .Q(currPixel[6])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i6.GSR = "DISABLED";
    FD1P3IX currPixel_679__i5 (.D(n37[5]), .SP(PIXEL_CLOCK_enable_25), .CD(n5345), 
            .CK(PIXEL_CLOCK), .Q(currPixel[5])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i5.GSR = "DISABLED";
    FD1P3IX currPixel_679__i4 (.D(n37[4]), .SP(PIXEL_CLOCK_enable_25), .CD(n5345), 
            .CK(PIXEL_CLOCK), .Q(currPixel[4])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i4.GSR = "DISABLED";
    FD1P3IX currPixel_679__i3 (.D(n37[3]), .SP(PIXEL_CLOCK_enable_25), .CD(n5345), 
            .CK(PIXEL_CLOCK), .Q(currPixel[3])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i3.GSR = "DISABLED";
    PFUMX i8380 (.BLUT(n11268), .ALUT(n11269), .C0(currBit[1]), .Z(n11272));
    FD1P3IX currPixel_679__i2 (.D(n37[2]), .SP(PIXEL_CLOCK_enable_25), .CD(n5345), 
            .CK(PIXEL_CLOCK), .Q(currPixel[2])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i2.GSR = "DISABLED";
    FD1P3IX currBit_680__i2 (.D(n21[2]), .SP(PIXEL_CLOCK_enable_13), .CD(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(currBit[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_680__i2.GSR = "DISABLED";
    FD1P3IX currBit_680__i1 (.D(n21[1]), .SP(PIXEL_CLOCK_enable_13), .CD(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(currBit[1]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_680__i1.GSR = "DISABLED";
    FD1P3IX currBit_680__i3 (.D(n21[3]), .SP(PIXEL_CLOCK_enable_13), .CD(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(currBit[3]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currBit_680__i3.GSR = "DISABLED";
    PFUMX i8381 (.BLUT(n11270), .ALUT(n11271), .C0(currBit[1]), .Z(n11273));
    FD1P3AX lastRow_i0_i0 (.D(MATRIX_CURRROW[0]), .SP(PIXEL_CLOCK_enable_20), 
            .CK(PIXEL_CLOCK), .Q(lastRow[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam lastRow_i0_i0.GSR = "DISABLED";
    PFUMX i8387 (.BLUT(n11275), .ALUT(n11276), .C0(currBit[1]), .Z(n11279));
    FD1S3AX currRow_i0_i0 (.D(n12[0]), .CK(PIXEL_CLOCK), .Q(MATRIX_CURRROW[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam currRow_i0_i0.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i1 (.D(n3), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5332), .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i1.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i4 (.D(n7), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i4.GSR = "DISABLED";
    FD1P3AY brightness_0__162 (.D(\BUS_data[0] ), .SP(LOGIC_CLOCK_N_116_enable_22), 
            .CK(LOGIC_CLOCK_N_116), .Q(\PWMArray[0][9] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam brightness_0__162.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i2 (.D(n3_adj_1219), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5332), .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i2.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i3 (.D(n13137), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i3.GSR = "DISABLED";
    FD1P3AY brightness_1__161 (.D(\BUS_data[1] ), .SP(LOGIC_CLOCK_N_116_enable_22), 
            .CK(LOGIC_CLOCK_N_116), .Q(\PWMArray[0][10] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam brightness_1__161.GSR = "DISABLED";
    FD1P3IX currPWMVal_i0_i5 (.D(n13138), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i5.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i12 (.D(currPWMVal_15__N_213[12]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i12.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i6 (.D(currPWMVal_15__N_213[6]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i6.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i3 (.D(n12333), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5332), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i3.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i6 (.D(n21[2]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i6.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i2 (.D(n21[1]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5332), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i2.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i5 (.D(n7_adj_1220), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i5.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i4 (.D(n7_adj_1221), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i4.GSR = "DISABLED";
    FD1P3IX currPWMCountMax__i7 (.D(currBit[2]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CD(n5322), .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i7.GSR = "DISABLED";
    CCU2D add_107_9 (.A0(currPWMCount[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9971), .COUT(n9972), .S0(currPWMCount_15__N_262[7]), 
          .S1(currPWMCount_15__N_262[8]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_9.INIT0 = 16'h5aaa;
    defparam add_107_9.INIT1 = 16'h5aaa;
    defparam add_107_9.INJECT1_0 = "NO";
    defparam add_107_9.INJECT1_1 = "NO";
    FD1P3AX MATRIX_ROWLAT_149 (.D(n12254), .SP(PIXEL_CLOCK_enable_15), .CK(PIXEL_CLOCK), 
            .Q(Matrix_LINE_SEL_Out_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam MATRIX_ROWLAT_149.GSR = "DISABLED";
    FD1P3BX currPWMCount_i15 (.D(currPWMCount_15__N_149[15]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i15.GSR = "DISABLED";
    FD1P3BX currPWMCount_i14 (.D(currPWMCount_15__N_149[14]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i14.GSR = "DISABLED";
    FD1P3BX currPWMCount_i13 (.D(currPWMCount_15__N_149[13]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i13.GSR = "DISABLED";
    FD1P3BX currPWMCount_i12 (.D(currPWMCount_15__N_149[12]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i12.GSR = "DISABLED";
    FD1P3BX currPWMCount_i11 (.D(currPWMCount_15__N_149[11]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i11.GSR = "DISABLED";
    FD1P3BX currPWMCount_i10 (.D(currPWMCount_15__N_149[10]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i10.GSR = "DISABLED";
    FD1P3BX currPWMCount_i9 (.D(currPWMCount_15__N_149[9]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i9.GSR = "DISABLED";
    FD1P3BX currPWMCount_i8 (.D(currPWMCount_15__N_149[8]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i8.GSR = "DISABLED";
    FD1P3BX currPWMCount_i7 (.D(currPWMCount_15__N_149[7]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i7.GSR = "DISABLED";
    FD1P3BX currPWMCount_i6 (.D(currPWMCount_15__N_149[6]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i6.GSR = "DISABLED";
    FD1P3BX currPWMCount_i5 (.D(currPWMCount_15__N_149[5]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i5.GSR = "DISABLED";
    FD1P3BX currPWMCount_i4 (.D(currPWMCount_15__N_149[4]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i4.GSR = "DISABLED";
    FD1P3BX currPWMCount_i3 (.D(currPWMCount_15__N_149[3]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i3.GSR = "DISABLED";
    FD1P3BX currPWMCount_i2 (.D(currPWMCount_15__N_149[2]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i2.GSR = "DISABLED";
    FD1P3BX currPWMCount_i1 (.D(currPWMCount_15__N_149[1]), .SP(LOGIC_CLOCK_enable_64), 
            .CK(LOGIC_CLOCK), .PD(Matrix_CTRL_Out_c_1), .Q(currPWMCount[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(202[3] 210[10])
    defparam currPWMCount_i1.GSR = "DISABLED";
    CCU2D add_7187_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n10116), 
          .S0(n1886));
    defparam add_7187_cout.INIT0 = 16'h0000;
    defparam add_7187_cout.INIT1 = 16'h0000;
    defparam add_7187_cout.INJECT1_0 = "NO";
    defparam add_7187_cout.INJECT1_1 = "NO";
    CCU2D add_7187_21 (.A0(\BUS_currGrantID[0] ), .B0(\BUS_currGrantID[1] ), 
          .C0(GND_net), .D0(GND_net), .A1(\BUS_currGrantID[0] ), .B1(\BUS_currGrantID[1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n10115), .COUT(n10116));
    defparam add_7187_21.INIT0 = 16'heeee;
    defparam add_7187_21.INIT1 = 16'heeee;
    defparam add_7187_21.INJECT1_0 = "NO";
    defparam add_7187_21.INJECT1_1 = "NO";
    PFUMX i8415 (.BLUT(n11303), .ALUT(n11304), .C0(currBit[1]), .Z(n11307));
    CCU2D add_7187_19 (.A0(n13158), .B0(n12344), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[18] ), 
          .D1(n12309), .CIN(n10114), .COUT(n10115));
    defparam add_7187_19.INIT0 = 16'h8888;
    defparam add_7187_19.INIT1 = 16'hff20;
    defparam add_7187_19.INJECT1_0 = "NO";
    defparam add_7187_19.INJECT1_1 = "NO";
    FD1P3AX currPWMCountMax__i13 (.D(currPWMCountMax_15__N_230[12]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i13.GSR = "DISABLED";
    CCU2D add_7187_17 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[15] ), .D0(n13150), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[16] ), .D1(n13151), 
          .CIN(n10113), .COUT(n10114));
    defparam add_7187_17.INIT0 = 16'h00ae;
    defparam add_7187_17.INIT1 = 16'h00ae;
    defparam add_7187_17.INJECT1_0 = "NO";
    defparam add_7187_17.INJECT1_1 = "NO";
    CCU2D sub_674_add_2_17 (.A0(currPWMCount[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10003), .S1(Matrix_CTRL_Out_c_2));
    defparam sub_674_add_2_17.INIT0 = 16'h5555;
    defparam sub_674_add_2_17.INIT1 = 16'h0000;
    defparam sub_674_add_2_17.INJECT1_0 = "NO";
    defparam sub_674_add_2_17.INJECT1_1 = "NO";
    FD1P3AX currPWMCountMax__i12 (.D(currPWMCountMax_15__N_230[11]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i12.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i11 (.D(currPWMCountMax_15__N_230[10]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i11.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i10 (.D(currPWMCountMax_15__N_230[9]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i10.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i9 (.D(currPWMCountMax_15__N_230[8]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i9.GSR = "DISABLED";
    FD1P3AX currPWMCountMax__i8 (.D(currPWMCountMax_15__N_230[7]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(\currPWMCountMax[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMCountMax__i8.GSR = "DISABLED";
    CCU2D add_7187_15 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[13] ), .D0(n13155), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[14] ), .D1(n13157), 
          .CIN(n10112), .COUT(n10113));
    defparam add_7187_15.INIT0 = 16'h00ae;
    defparam add_7187_15.INIT1 = 16'h00ae;
    defparam add_7187_15.INJECT1_0 = "NO";
    defparam add_7187_15.INJECT1_1 = "NO";
    FD1P3AX currPWMVal_i0_i11 (.D(currPWMVal_15__N_213[11]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i11.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i10 (.D(currPWMVal_15__N_213[10]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i10.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i9 (.D(currPWMVal_15__N_213[9]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i9.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i8 (.D(currPWMVal_15__N_213[8]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i8.GSR = "DISABLED";
    FD1P3AX currPWMVal_i0_i7 (.D(currPWMVal_15__N_213[7]), .SP(PIXEL_CLOCK_N_302_enable_26), 
            .CK(PIXEL_CLOCK_N_302), .Q(currPWMVal[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(188[3] 194[10])
    defparam currPWMVal_i0_i7.GSR = "DISABLED";
    CCU2D sub_674_add_2_15 (.A0(currPWMCount[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10002), .COUT(n10003));
    defparam sub_674_add_2_15.INIT0 = 16'h5555;
    defparam sub_674_add_2_15.INIT1 = 16'h5555;
    defparam sub_674_add_2_15.INJECT1_0 = "NO";
    defparam sub_674_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_674_add_2_13 (.A0(currPWMCount[11]), .B0(currPWMVal[11]), 
          .C0(GND_net), .D0(GND_net), .A1(currPWMCount[12]), .B1(currPWMVal[12]), 
          .C1(GND_net), .D1(GND_net), .CIN(n10001), .COUT(n10002));
    defparam sub_674_add_2_13.INIT0 = 16'h5999;
    defparam sub_674_add_2_13.INIT1 = 16'h5999;
    defparam sub_674_add_2_13.INJECT1_0 = "NO";
    defparam sub_674_add_2_13.INJECT1_1 = "NO";
    CCU2D add_7187_13 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[11] ), .D0(n13156), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[12] ), .D1(n13142), 
          .CIN(n10111), .COUT(n10112));
    defparam add_7187_13.INIT0 = 16'h00ae;
    defparam add_7187_13.INIT1 = 16'h00ae;
    defparam add_7187_13.INJECT1_0 = "NO";
    defparam add_7187_13.INJECT1_1 = "NO";
    CCU2D sub_674_add_2_11 (.A0(currPWMCount[9]), .B0(currPWMVal[9]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[10]), .B1(currPWMVal[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n10000), .COUT(n10001));
    defparam sub_674_add_2_11.INIT0 = 16'h5999;
    defparam sub_674_add_2_11.INIT1 = 16'h5999;
    defparam sub_674_add_2_11.INJECT1_0 = "NO";
    defparam sub_674_add_2_11.INJECT1_1 = "NO";
    PFUMX i8388 (.BLUT(n11277), .ALUT(n11278), .C0(currBit[1]), .Z(n11280));
    CCU2D add_7187_11 (.A0(\BUS_ADDR_INTERNAL[9] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13144), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[10] ), .D1(n13143), 
          .CIN(n10110), .COUT(n10111));
    defparam add_7187_11.INIT0 = 16'h00dc;
    defparam add_7187_11.INIT1 = 16'hff51;
    defparam add_7187_11.INJECT1_0 = "NO";
    defparam add_7187_11.INJECT1_1 = "NO";
    CCU2D sub_674_add_2_9 (.A0(currPWMCount[7]), .B0(currPWMVal[7]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[8]), .B1(currPWMVal[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9999), .COUT(n10000));
    defparam sub_674_add_2_9.INIT0 = 16'h5999;
    defparam sub_674_add_2_9.INIT1 = 16'h5999;
    defparam sub_674_add_2_9.INJECT1_0 = "NO";
    defparam sub_674_add_2_9.INJECT1_1 = "NO";
    CCU2D add_7187_9 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[7] ), .D0(n13147), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[8] ), .D1(n13154), 
          .CIN(n10109), .COUT(n10110));
    defparam add_7187_9.INIT0 = 16'hff51;
    defparam add_7187_9.INIT1 = 16'h00ae;
    defparam add_7187_9.INJECT1_0 = "NO";
    defparam add_7187_9.INJECT1_1 = "NO";
    LUT4 i14_4_lut (.A(currPWMCount[10]), .B(n28), .C(n22_adj_1222), .D(currPWMCount[12]), 
         .Z(n30)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i14_4_lut.init = 16'h8000;
    CCU2D add_7187_7 (.A0(\BUS_ADDR_INTERNAL[5] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13145), .A1(\BUS_currGrantID[1] ), 
          .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[6] ), .D1(n13146), 
          .CIN(n10108), .COUT(n10109));
    defparam add_7187_7.INIT0 = 16'h00dc;
    defparam add_7187_7.INIT1 = 16'h00ae;
    defparam add_7187_7.INJECT1_0 = "NO";
    defparam add_7187_7.INJECT1_1 = "NO";
    CCU2D add_7187_5 (.A0(\BUS_currGrantID[1] ), .B0(\BUS_currGrantID[0] ), 
          .C0(\BUS_ADDR_INTERNAL[3] ), .D0(n13148), .A1(\BUS_ADDR_INTERNAL[4] ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13153), 
          .CIN(n10107), .COUT(n10108));
    defparam add_7187_5.INIT0 = 16'h00ae;
    defparam add_7187_5.INIT1 = 16'h00dc;
    defparam add_7187_5.INJECT1_0 = "NO";
    defparam add_7187_5.INJECT1_1 = "NO";
    PFUMX i8394 (.BLUT(n11282), .ALUT(n11283), .C0(currBit[1]), .Z(n11286));
    CCU2D add_7187_3 (.A0(\BUS_ADDR_INTERNAL[1] ), .B0(\BUS_currGrantID[1] ), 
          .C0(\BUS_currGrantID[0] ), .D0(n13149), .A1(\BUS_ADDR_INTERNAL[2] ), 
          .B1(\BUS_currGrantID[1] ), .C1(\BUS_currGrantID[0] ), .D1(n13152), 
          .CIN(n10106), .COUT(n10107));
    defparam add_7187_3.INIT0 = 16'h00dc;
    defparam add_7187_3.INIT1 = 16'h00dc;
    defparam add_7187_3.INJECT1_0 = "NO";
    defparam add_7187_3.INJECT1_1 = "NO";
    CCU2D add_7187_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\BUS_currGrantID[1] ), .B1(\BUS_currGrantID[0] ), .C1(\BUS_ADDR_INTERNAL[0] ), 
          .D1(n12299), .COUT(n10106));
    defparam add_7187_1.INIT0 = 16'hF000;
    defparam add_7187_1.INIT1 = 16'h00ae;
    defparam add_7187_1.INJECT1_0 = "NO";
    defparam add_7187_1.INJECT1_1 = "NO";
    FD1P3AX currPixel_679__i0 (.D(n47[0]), .SP(PIXEL_CLOCK_enable_25), .CK(PIXEL_CLOCK), 
            .Q(currPixel[0])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i0.GSR = "DISABLED";
    CCU2D sub_674_add_2_7 (.A0(currPWMCount[5]), .B0(currPWMVal[5]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[6]), .B1(currPWMVal[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9998), .COUT(n9999));
    defparam sub_674_add_2_7.INIT0 = 16'h5999;
    defparam sub_674_add_2_7.INIT1 = 16'h5999;
    defparam sub_674_add_2_7.INJECT1_0 = "NO";
    defparam sub_674_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_674_add_2_5 (.A0(currPWMCount[3]), .B0(currPWMVal[3]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[4]), .B1(currPWMVal[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9997), .COUT(n9998));
    defparam sub_674_add_2_5.INIT0 = 16'h5999;
    defparam sub_674_add_2_5.INIT1 = 16'h5999;
    defparam sub_674_add_2_5.INJECT1_0 = "NO";
    defparam sub_674_add_2_5.INJECT1_1 = "NO";
    PFUMX i8395 (.BLUT(n11284), .ALUT(n11285), .C0(currBit[1]), .Z(n11287));
    PFUMX i8401 (.BLUT(n11289), .ALUT(n11290), .C0(currBit[1]), .Z(n11293));
    PFUMX i8402 (.BLUT(n11291), .ALUT(n11292), .C0(currBit[1]), .Z(n11294));
    CCU2D sub_674_add_2_3 (.A0(currPWMCount[1]), .B0(currPWMVal[1]), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[2]), .B1(currPWMVal[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n9996), .COUT(n9997));
    defparam sub_674_add_2_3.INIT0 = 16'h5999;
    defparam sub_674_add_2_3.INIT1 = 16'h5999;
    defparam sub_674_add_2_3.INJECT1_0 = "NO";
    defparam sub_674_add_2_3.INJECT1_1 = "NO";
    PFUMX i8408 (.BLUT(n11296), .ALUT(n11297), .C0(currBit[1]), .Z(n11300));
    PFUMX i8409 (.BLUT(n11298), .ALUT(n11299), .C0(currBit[1]), .Z(n11301));
    CCU2D sub_674_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(currPWMCount[0]), .B1(currPWMVal[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n9996));
    defparam sub_674_add_2_1.INIT0 = 16'h0000;
    defparam sub_674_add_2_1.INIT1 = 16'h5999;
    defparam sub_674_add_2_1.INJECT1_0 = "NO";
    defparam sub_674_add_2_1.INJECT1_1 = "NO";
    LUT4 i1024_1_lut (.A(MATRIX_CURRROW[0]), .Z(currReadRow[0])) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1024_1_lut.init = 16'h5555;
    LUT4 i8407_3_lut (.A(\RED[1] [6]), .B(\RED[1] [7]), .C(currBit[0]), 
         .Z(n11299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8407_3_lut.init = 16'hcaca;
    LUT4 mux_92_Mux_7_i15_4_lut_4_lut (.A(currBit[0]), .B(currBit[1]), .C(currBit[2]), 
         .D(currBit[3]), .Z(currPWMCountMax_15__N_230[7])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B (C+!(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(191[36:65])
    defparam mux_92_Mux_7_i15_4_lut_4_lut.init = 16'h01e0;
    LUT4 i180_4_lut (.A(n12260), .B(currPixel[7]), .C(n12231), .D(n12249), 
         .Z(n1095)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C+(D))+!B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(147[4] 185[11])
    defparam i180_4_lut.init = 16'h880c;
    LUT4 currBit_3__I_0_164_i15_4_lut (.A(n11246), .B(n8), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_11)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(137[26:55])
    defparam currBit_3__I_0_164_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_164_i8_3_lut (.A(\BLUE[3] [8]), .B(\BLUE[3] [9]), 
         .C(currBit[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(137[26:55])
    defparam currBit_3__I_0_164_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_165_i15_4_lut (.A(n11253), .B(n8_adj_1223), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_10)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(136[27:56])
    defparam currBit_3__I_0_165_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_165_i8_3_lut (.A(\GREEN[3] [8]), .B(\GREEN[3] [9]), 
         .C(currBit[0]), .Z(n8_adj_1223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(136[27:56])
    defparam currBit_3__I_0_165_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_166_i15_4_lut (.A(n11260), .B(n8_adj_1224), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_9)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(135[24:53])
    defparam currBit_3__I_0_166_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_166_i8_3_lut (.A(\RED[3] [8]), .B(\RED[3] [9]), 
         .C(currBit[0]), .Z(n8_adj_1224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(135[24:53])
    defparam currBit_3__I_0_166_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_167_i15_4_lut (.A(n11267), .B(n8_adj_1225), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_8)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(133[25:54])
    defparam currBit_3__I_0_167_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_167_i8_3_lut (.A(\BLUE[2] [8]), .B(\BLUE[2] [9]), 
         .C(currBit[0]), .Z(n8_adj_1225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(133[25:54])
    defparam currBit_3__I_0_167_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_168_i15_4_lut (.A(n11274), .B(n8_adj_1226), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_7)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(132[26:55])
    defparam currBit_3__I_0_168_i15_4_lut.init = 16'hca0a;
    LUT4 i4_4_lut (.A(currPixel[4]), .B(currPixel[5]), .C(currPixel[2]), 
         .D(currPixel[6]), .Z(n10_adj_1227)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 currBit_3__I_0_168_i8_3_lut (.A(\GREEN[2] [8]), .B(\GREEN[2] [9]), 
         .C(currBit[0]), .Z(n8_adj_1226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(132[26:55])
    defparam currBit_3__I_0_168_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_169_i15_4_lut (.A(n11281), .B(n8_adj_1228), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_6)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(131[24:53])
    defparam currBit_3__I_0_169_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_169_i8_3_lut (.A(\RED[2] [8]), .B(\RED[2] [9]), 
         .C(currBit[0]), .Z(n8_adj_1228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(131[24:53])
    defparam currBit_3__I_0_169_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_170_i15_4_lut (.A(n11288), .B(n8_adj_1229), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_5)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(129[25:54])
    defparam currBit_3__I_0_170_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_170_i8_3_lut (.A(\BLUE[1] [8]), .B(\BLUE[1] [9]), 
         .C(currBit[0]), .Z(n8_adj_1229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(129[25:54])
    defparam currBit_3__I_0_170_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_171_i15_4_lut (.A(n11295), .B(n8_adj_1230), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_4)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(128[26:55])
    defparam currBit_3__I_0_171_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_2__bdd_4_lut_9524 (.A(currBit[2]), .B(n12306), .C(n14), 
         .D(currBit[3]), .Z(currPWMVal_15__N_213[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam currBit_2__bdd_4_lut_9524.init = 16'hf088;
    LUT4 currBit_3__I_0_171_i8_3_lut (.A(\GREEN[1] [8]), .B(\GREEN[1] [9]), 
         .C(currBit[0]), .Z(n8_adj_1230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(128[26:55])
    defparam currBit_3__I_0_171_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_172_i15_4_lut (.A(n11302), .B(n8_adj_1231), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_3)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(127[24:53])
    defparam currBit_3__I_0_172_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_172_i8_3_lut (.A(\RED[1] [8]), .B(\RED[1] [9]), 
         .C(currBit[0]), .Z(n8_adj_1231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(127[24:53])
    defparam currBit_3__I_0_172_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_173_i15_4_lut (.A(n11309), .B(n8_adj_1232), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_2)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(125[25:54])
    defparam currBit_3__I_0_173_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_173_i8_3_lut (.A(\BLUE[0] [8]), .B(\BLUE[0] [9]), 
         .C(currBit[0]), .Z(n8_adj_1232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(125[25:54])
    defparam currBit_3__I_0_173_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_174_i15_4_lut (.A(n11316), .B(n8_adj_1233), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_1)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(124[26:55])
    defparam currBit_3__I_0_174_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_174_i8_3_lut (.A(\GREEN[0] [8]), .B(\GREEN[0] [9]), 
         .C(currBit[0]), .Z(n8_adj_1233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(124[26:55])
    defparam currBit_3__I_0_174_i8_3_lut.init = 16'hcaca;
    LUT4 currBit_3__I_0_184_i15_4_lut (.A(n11323), .B(n8_adj_1234), .C(currBit[3]), 
         .D(n12349), .Z(Matrix_DATA_Out_c_0)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(123[24:53])
    defparam currBit_3__I_0_184_i15_4_lut.init = 16'hca0a;
    LUT4 currBit_3__I_0_184_i8_3_lut (.A(\RED[0] [8]), .B(\RED[0] [9]), 
         .C(currBit[0]), .Z(n8_adj_1234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(123[24:53])
    defparam currBit_3__I_0_184_i8_3_lut.init = 16'hcaca;
    LUT4 i8635_4_lut (.A(MATRIX_CURRROW[3]), .B(MATRIX_CURRROW[2]), .C(MATRIX_CURRROW[0]), 
         .D(n6), .Z(Matrix_LINE_SEL_Out_c_2)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(141[29:46])
    defparam i8635_4_lut.init = 16'h0001;
    LUT4 i1_2_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[4]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(141[29:46])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i4566_2_lut (.A(PIXEL_CLOCK), .B(MATRIX_CLKEN_LAT), .Z(Matrix_CTRL_Out_c_0)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(197[18:66])
    defparam i4566_2_lut.init = 16'h8888;
    LUT4 i8428_3_lut (.A(\RED[0] [6]), .B(\RED[0] [7]), .C(currBit[0]), 
         .Z(n11320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8428_3_lut.init = 16'hcaca;
    LUT4 i8427_3_lut (.A(\RED[0] [4]), .B(\RED[0] [5]), .C(currBit[0]), 
         .Z(n11319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8427_3_lut.init = 16'hcaca;
    LUT4 i8426_3_lut (.A(\RED[0] [2]), .B(\RED[0] [3]), .C(currBit[0]), 
         .Z(n11318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8426_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(MATRIX_CURRROW[3]), .B(n12311), .C(MATRIX_CURRROW[4]), 
         .D(\lastReadRow[4] ), .Z(n10349)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i2_3_lut_4_lut.init = 16'h8778;
    LUT4 n8_bdd_4_lut (.A(n12336), .B(currBit[3]), .C(\PWMArray[0][10] ), 
         .D(currBit[0]), .Z(n12135)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B+((D)+!C))) */ ;
    defparam n8_bdd_4_lut.init = 16'h88b8;
    LUT4 i8425_3_lut (.A(\RED[0] [0]), .B(\RED[0] [1]), .C(currBit[0]), 
         .Z(n11317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8425_3_lut.init = 16'hcaca;
    LUT4 i8421_3_lut (.A(\GREEN[0] [6]), .B(\GREEN[0] [7]), .C(currBit[0]), 
         .Z(n11313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8421_3_lut.init = 16'hcaca;
    LUT4 BUS_VALID_I_7_2_lut_rep_195 (.A(BUS_VALID_N_113), .B(n1886), .Z(n12221)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(261[29:83])
    defparam BUS_VALID_I_7_2_lut_rep_195.init = 16'h2222;
    LUT4 i8590_2_lut_3_lut_4_lut (.A(BUS_VALID_N_113), .B(n1886), .C(n13141), 
         .D(n87), .Z(LOGIC_CLOCK_N_116_enable_22)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(261[29:83])
    defparam i8590_2_lut_3_lut_4_lut.init = 16'h0020;
    CCU2D currPixel_679_add_4_9 (.A0(currPixel[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n10037), .S0(n37[7]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679_add_4_9.INIT0 = 16'hfaaa;
    defparam currPixel_679_add_4_9.INIT1 = 16'h0000;
    defparam currPixel_679_add_4_9.INJECT1_0 = "NO";
    defparam currPixel_679_add_4_9.INJECT1_1 = "NO";
    LUT4 i8406_3_lut (.A(\RED[1] [4]), .B(\RED[1] [5]), .C(currBit[0]), 
         .Z(n11298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8406_3_lut.init = 16'hcaca;
    LUT4 i8420_3_lut (.A(\GREEN[0] [4]), .B(\GREEN[0] [5]), .C(currBit[0]), 
         .Z(n11312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8420_3_lut.init = 16'hcaca;
    LUT4 i8419_3_lut (.A(\GREEN[0] [2]), .B(\GREEN[0] [3]), .C(currBit[0]), 
         .Z(n11311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8419_3_lut.init = 16'hcaca;
    LUT4 i8418_3_lut (.A(\GREEN[0] [0]), .B(\GREEN[0] [1]), .C(currBit[0]), 
         .Z(n11310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8418_3_lut.init = 16'hcaca;
    CCU2D currPixel_679_add_4_7 (.A0(currPixel[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10036), .COUT(n10037), .S0(n37[5]), .S1(n37[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679_add_4_7.INIT0 = 16'hfaaa;
    defparam currPixel_679_add_4_7.INIT1 = 16'hfaaa;
    defparam currPixel_679_add_4_7.INJECT1_0 = "NO";
    defparam currPixel_679_add_4_7.INJECT1_1 = "NO";
    CCU2D add_107_7 (.A0(currPWMCount[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9970), .COUT(n9971), .S0(currPWMCount_15__N_262[5]), 
          .S1(currPWMCount_15__N_262[6]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_7.INIT0 = 16'h5aaa;
    defparam add_107_7.INIT1 = 16'h5aaa;
    defparam add_107_7.INJECT1_0 = "NO";
    defparam add_107_7.INJECT1_1 = "NO";
    LUT4 currBit_2__bdd_4_lut_9635 (.A(currBit[2]), .B(n12334), .C(n12359), 
         .D(currBit[1]), .Z(n13137)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam currBit_2__bdd_4_lut_9635.init = 16'h44f0;
    LUT4 currBit_2__bdd_4_lut (.A(currBit[2]), .B(n12334), .C(n12357), 
         .D(currBit[1]), .Z(n13138)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam currBit_2__bdd_4_lut.init = 16'hf088;
    CCU2D currPixel_679_add_4_5 (.A0(currPixel[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10035), .COUT(n10036), .S0(n37[3]), .S1(n37[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679_add_4_5.INIT0 = 16'hfaaa;
    defparam currPixel_679_add_4_5.INIT1 = 16'hfaaa;
    defparam currPixel_679_add_4_5.INJECT1_0 = "NO";
    defparam currPixel_679_add_4_5.INJECT1_1 = "NO";
    CCU2D currPixel_679_add_4_3 (.A0(currPixel[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n10034), .COUT(n10035), .S0(n37[1]), .S1(n37[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679_add_4_3.INIT0 = 16'hfaaa;
    defparam currPixel_679_add_4_3.INIT1 = 16'hfaaa;
    defparam currPixel_679_add_4_3.INJECT1_0 = "NO";
    defparam currPixel_679_add_4_3.INJECT1_1 = "NO";
    FD1P3AX lastRow_i0_i1 (.D(MATRIX_CURRROW[1]), .SP(PIXEL_CLOCK_enable_20), 
            .CK(PIXEL_CLOCK), .Q(lastRow[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam lastRow_i0_i1.GSR = "DISABLED";
    FD1P3AX lastRow_i0_i2 (.D(MATRIX_CURRROW[2]), .SP(PIXEL_CLOCK_enable_20), 
            .CK(PIXEL_CLOCK), .Q(lastRow[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam lastRow_i0_i2.GSR = "DISABLED";
    FD1P3AX lastRow_i0_i3 (.D(MATRIX_CURRROW[3]), .SP(PIXEL_CLOCK_enable_20), 
            .CK(PIXEL_CLOCK), .Q(lastRow[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam lastRow_i0_i3.GSR = "DISABLED";
    FD1P3AX lastRow_i0_i4 (.D(MATRIX_CURRROW[4]), .SP(PIXEL_CLOCK_enable_20), 
            .CK(PIXEL_CLOCK), .Q(lastRow[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam lastRow_i0_i4.GSR = "DISABLED";
    FD1P3AX currRow_i0_i1 (.D(currReadRow[1]), .SP(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(MATRIX_CURRROW[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam currRow_i0_i1.GSR = "DISABLED";
    FD1P3AX currRow_i0_i2 (.D(currReadRow[2]), .SP(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(MATRIX_CURRROW[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam currRow_i0_i2.GSR = "DISABLED";
    FD1P3AX currRow_i0_i3 (.D(currReadRow[3]), .SP(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(MATRIX_CURRROW[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam currRow_i0_i3.GSR = "DISABLED";
    FD1P3AX currRow_i0_i4 (.D(currReadRow[4]), .SP(PIXEL_CLOCK_enable_24), 
            .CK(PIXEL_CLOCK), .Q(MATRIX_CURRROW[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam currRow_i0_i4.GSR = "DISABLED";
    FD1S3AX currPixel_679__i1 (.D(n12047), .CK(PIXEL_CLOCK), .Q(currPixel[1])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i1.GSR = "DISABLED";
    CCU2D add_107_5 (.A0(currPWMCount[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9969), .COUT(n9970), .S0(currPWMCount_15__N_262[3]), 
          .S1(currPWMCount_15__N_262[4]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_5.INIT0 = 16'h5aaa;
    defparam add_107_5.INIT1 = 16'h5aaa;
    defparam add_107_5.INJECT1_0 = "NO";
    defparam add_107_5.INJECT1_1 = "NO";
    CCU2D currPixel_679_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPixel[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n10034), .S1(n37[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679_add_4_1.INIT0 = 16'hF000;
    defparam currPixel_679_add_4_1.INIT1 = 16'h0555;
    defparam currPixel_679_add_4_1.INJECT1_0 = "NO";
    defparam currPixel_679_add_4_1.INJECT1_1 = "NO";
    LUT4 i8627_2_lut_rep_229_3_lut (.A(currPixel[0]), .B(n12330), .C(currPixel[1]), 
         .Z(PIXEL_CLOCK_N_302_enable_26)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i8627_2_lut_rep_229_3_lut.init = 16'h2020;
    LUT4 i2734_2_lut_3_lut_4_lut (.A(currPixel[0]), .B(n12330), .C(currBit[3]), 
         .D(currPixel[1]), .Z(n5322)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i2734_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_234_3_lut (.A(currPixel[0]), .B(n12330), .C(currPixel[1]), 
         .Z(n12260)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i1_2_lut_rep_234_3_lut.init = 16'hfdfd;
    LUT4 i8720_2_lut_2_lut_3_lut_4_lut (.A(currPixel[1]), .B(n12275), .C(n12231), 
         .D(currPixel[7]), .Z(PIXEL_CLOCK_enable_25)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(150[10:27])
    defparam i8720_2_lut_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i8578_2_lut_3_lut_4_lut (.A(currPixel[0]), .B(n12330), .C(currBit[0]), 
         .D(currPixel[1]), .Z(n7141)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i8578_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_217_3_lut_4_lut (.A(currPixel[0]), .B(n12330), .C(MATRIX_ROWCLK_N_289), 
         .D(currPixel[1]), .Z(n12243)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i1_2_lut_rep_217_3_lut_4_lut.init = 16'h0020;
    LUT4 i8414_3_lut (.A(\BLUE[0] [6]), .B(\BLUE[0] [7]), .C(currBit[0]), 
         .Z(n11306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8414_3_lut.init = 16'hcaca;
    LUT4 i8413_3_lut (.A(\BLUE[0] [4]), .B(\BLUE[0] [5]), .C(currBit[0]), 
         .Z(n11305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8413_3_lut.init = 16'hcaca;
    PFUMX i8416 (.BLUT(n11305), .ALUT(n11306), .C0(currBit[1]), .Z(n11308));
    LUT4 i8412_3_lut (.A(\BLUE[0] [2]), .B(\BLUE[0] [3]), .C(currBit[0]), 
         .Z(n11304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8412_3_lut.init = 16'hcaca;
    LUT4 mux_91_Mux_5_i7_3_lut_4_lut_then_4_lut (.A(currBit[2]), .B(\PWMArray[0][9] ), 
         .C(currBit[0]), .D(\PWMArray[0][12] ), .Z(n12357)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam mux_91_Mux_5_i7_3_lut_4_lut_then_4_lut.init = 16'h5808;
    LUT4 i8411_3_lut (.A(\BLUE[0] [0]), .B(\BLUE[0] [1]), .C(currBit[0]), 
         .Z(n11303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8411_3_lut.init = 16'hcaca;
    LUT4 i1026_2_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), .Z(currReadRow[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1026_2_lut.init = 16'h6666;
    LUT4 VRAM_READ_ADDR_7__I_0_1_lut (.A(VRAM_READ_ADDR[7]), .Z(VRAM_WRITE_ADDR[7])) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(236[24:44])
    defparam VRAM_READ_ADDR_7__I_0_1_lut.init = 16'h5555;
    LUT4 mux_91_Mux_3_i7_3_lut_4_lut_else_2_lut (.A(currBit[2]), .B(\PWMArray[0][12] ), 
         .C(currBit[0]), .D(\PWMArray[0][9] ), .Z(n12359)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)))) */ ;
    defparam mux_91_Mux_3_i7_3_lut_4_lut_else_2_lut.init = 16'h4a40;
    LUT4 mux_91_Mux_9_i7_3_lut_4_lut_4_lut (.A(currBit[1]), .B(n12335), 
         .C(currBit[2]), .D(n12340), .Z(n7_adj_1235)) /* synthesis lut_function=(A (B (C))+!A !(C+!(D))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(273[3] 280[10])
    defparam mux_91_Mux_9_i7_3_lut_4_lut_4_lut.init = 16'h8580;
    LUT4 i4829_2_lut_4_lut (.A(n12335), .B(n12334), .C(currBit[1]), .D(currBit[2]), 
         .Z(n7_adj_1236)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i4829_2_lut_4_lut.init = 16'hca00;
    FD1P3AX currPixel_679__i7 (.D(n47[7]), .SP(PIXEL_CLOCK_enable_25), .CK(PIXEL_CLOCK), 
            .Q(currPixel[7])) /* synthesis syn_use_carry_chain=1 */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam currPixel_679__i7.GSR = "DISABLED";
    LUT4 mux_91_Mux_4_i7_4_lut_4_lut (.A(n12336), .B(currBit[1]), .C(currBit[2]), 
         .D(n12337), .Z(n7)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B+!(C (D))))) */ ;
    defparam mux_91_Mux_4_i7_4_lut_4_lut.init = 16'h3808;
    LUT4 currPixel_679_mux_6_i1_3_lut_4_lut (.A(currPixel[1]), .B(n12275), 
         .C(n1095), .D(n37[0]), .Z(n47[0])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam currPixel_679_mux_6_i1_3_lut_4_lut.init = 16'h2f20;
    LUT4 currPixel_679_mux_6_i8_3_lut_4_lut (.A(currPixel[1]), .B(n12275), 
         .C(n1095), .D(n37[7]), .Z(n47[7])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam currPixel_679_mux_6_i8_3_lut_4_lut.init = 16'h2f20;
    LUT4 i8405_3_lut (.A(\RED[1] [2]), .B(\RED[1] [3]), .C(currBit[0]), 
         .Z(n11297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8405_3_lut.init = 16'hcaca;
    PFUMX i8422 (.BLUT(n11310), .ALUT(n11311), .C0(currBit[1]), .Z(n11314));
    LUT4 i8404_3_lut (.A(\RED[1] [0]), .B(\RED[1] [1]), .C(currBit[0]), 
         .Z(n11296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8404_3_lut.init = 16'hcaca;
    LUT4 i8400_3_lut (.A(\GREEN[1] [6]), .B(\GREEN[1] [7]), .C(currBit[0]), 
         .Z(n11292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8400_3_lut.init = 16'hcaca;
    LUT4 i8399_3_lut (.A(\GREEN[1] [4]), .B(\GREEN[1] [5]), .C(currBit[0]), 
         .Z(n11291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8399_3_lut.init = 16'hcaca;
    LUT4 i8718_4_lut_4_lut (.A(n12231), .B(n26), .C(n30), .D(n25), .Z(LOGIC_CLOCK_enable_64)) /* synthesis lut_function=((B (C (D)))+!A) */ ;
    defparam i8718_4_lut_4_lut.init = 16'hd555;
    LUT4 i8398_3_lut (.A(\GREEN[1] [2]), .B(\GREEN[1] [3]), .C(currBit[0]), 
         .Z(n11290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8398_3_lut.init = 16'hcaca;
    LUT4 i8397_3_lut (.A(\GREEN[1] [0]), .B(\GREEN[1] [1]), .C(currBit[0]), 
         .Z(n11289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8397_3_lut.init = 16'hcaca;
    LUT4 i8393_3_lut (.A(\BLUE[1] [6]), .B(\BLUE[1] [7]), .C(currBit[0]), 
         .Z(n11285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8393_3_lut.init = 16'hcaca;
    LUT4 i8392_3_lut (.A(\BLUE[1] [4]), .B(\BLUE[1] [5]), .C(currBit[0]), 
         .Z(n11284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8392_3_lut.init = 16'hcaca;
    LUT4 i2736_3_lut_4_lut (.A(currPixel[1]), .B(n12285), .C(currBit[3]), 
         .D(currBit[2]), .Z(n5332)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i2736_3_lut_4_lut.init = 16'h2220;
    LUT4 i8391_3_lut (.A(\BLUE[1] [2]), .B(\BLUE[1] [3]), .C(currBit[0]), 
         .Z(n11283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8391_3_lut.init = 16'hcaca;
    LUT4 i8390_3_lut (.A(\BLUE[1] [0]), .B(\BLUE[1] [1]), .C(currBit[0]), 
         .Z(n11282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8390_3_lut.init = 16'hcaca;
    LUT4 i8716_2_lut_rep_323 (.A(currBit[1]), .B(currBit[2]), .Z(n12349)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i8716_2_lut_rep_323.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(\PWMArray[0][9] ), 
         .D(currBit[0]), .Z(n14_adj_1237)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i789_2_lut_rep_255_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), 
         .C(currBit[3]), .D(currBit[0]), .Z(n12281)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i789_2_lut_rep_255_3_lut_4_lut.init = 16'hf0e0;
    LUT4 LED_c_bdd_2_lut_3_lut (.A(currBit[1]), .B(currBit[2]), .C(n12135), 
         .Z(currPWMVal_15__N_213[10])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam LED_c_bdd_2_lut_3_lut.init = 16'h1010;
    LUT4 i8386_3_lut (.A(\RED[2] [6]), .B(\RED[2] [7]), .C(currBit[0]), 
         .Z(n11278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8386_3_lut.init = 16'hcaca;
    LUT4 LED_c_bdd_2_lut_8771_3_lut (.A(currBit[1]), .B(currBit[2]), .C(n11718), 
         .Z(currPWMVal_15__N_213[11])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam LED_c_bdd_2_lut_8771_3_lut.init = 16'h1010;
    LUT4 i4_4_lut_adj_121 (.A(n7_adj_1238), .B(lastRow[2]), .C(n6_adj_1239), 
         .D(MATRIX_CURRROW[2]), .Z(MATRIX_ROWCLK_N_289)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(160[13:30])
    defparam i4_4_lut_adj_121.init = 16'hfbfe;
    LUT4 i2_4_lut (.A(lastRow[3]), .B(lastRow[0]), .C(MATRIX_CURRROW[3]), 
         .D(MATRIX_CURRROW[0]), .Z(n7_adj_1238)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(160[13:30])
    defparam i2_4_lut.init = 16'h7bde;
    LUT4 i1_4_lut (.A(lastRow[1]), .B(lastRow[4]), .C(MATRIX_CURRROW[1]), 
         .D(MATRIX_CURRROW[4]), .Z(n6_adj_1239)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(160[13:30])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i8575_2_lut_rep_272_3_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .Z(n12298)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i8575_2_lut_rep_272_3_lut.init = 16'h0101;
    LUT4 i8385_3_lut (.A(\RED[2] [4]), .B(\RED[2] [5]), .C(currBit[0]), 
         .Z(n11277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8385_3_lut.init = 16'hcaca;
    LUT4 i8384_3_lut (.A(\RED[2] [2]), .B(\RED[2] [3]), .C(currBit[0]), 
         .Z(n11276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8384_3_lut.init = 16'hcaca;
    LUT4 i4880_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .D(currBit[0]), .Z(currPWMCountMax_15__N_230[11])) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;
    defparam i4880_3_lut_4_lut.init = 16'h1001;
    LUT4 i8624_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[0]), 
         .D(currBit[3]), .Z(currPWMCountMax_15__N_230[10])) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i8624_3_lut_4_lut.init = 16'h1101;
    LUT4 i2_4_lut_adj_122 (.A(MATRIX_CURRROW[2]), .B(\lastReadRow[3] ), 
         .C(n12342), .D(MATRIX_CURRROW[3]), .Z(n10350)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i2_4_lut_adj_122.init = 16'h936c;
    LUT4 mux_92_Mux_8_i15_4_lut_3_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[3]), 
         .Z(currPWMCountMax_15__N_230[8])) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_92_Mux_8_i15_4_lut_3_lut.init = 16'h1818;
    LUT4 i8383_3_lut (.A(\RED[2] [0]), .B(\RED[2] [1]), .C(currBit[0]), 
         .Z(n11275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8383_3_lut.init = 16'hcaca;
    LUT4 i8379_3_lut (.A(\GREEN[2] [6]), .B(\GREEN[2] [7]), .C(currBit[0]), 
         .Z(n11271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8379_3_lut.init = 16'hcaca;
    LUT4 i8378_3_lut (.A(\GREEN[2] [4]), .B(\GREEN[2] [5]), .C(currBit[0]), 
         .Z(n11270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8378_3_lut.init = 16'hcaca;
    LUT4 i8377_3_lut (.A(\GREEN[2] [2]), .B(\GREEN[2] [3]), .C(currBit[0]), 
         .Z(n11269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8377_3_lut.init = 16'hcaca;
    LUT4 i8376_3_lut (.A(\GREEN[2] [0]), .B(\GREEN[2] [1]), .C(currBit[0]), 
         .Z(n11268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8376_3_lut.init = 16'hcaca;
    CCU2D add_107_17 (.A0(currPWMCount[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n9975), .S0(currPWMCount_15__N_262[15]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_17.INIT0 = 16'h5aaa;
    defparam add_107_17.INIT1 = 16'h0000;
    defparam add_107_17.INJECT1_0 = "NO";
    defparam add_107_17.INJECT1_1 = "NO";
    LUT4 i7202_2_lut (.A(currBit[1]), .B(currBit[0]), .Z(n21[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i7202_2_lut.init = 16'h6666;
    LUT4 i1102_1_lut (.A(currPixel[1]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam i1102_1_lut.init = 16'h5555;
    LUT4 i8724_2_lut_3_lut_4_lut (.A(currBit[1]), .B(currBit[2]), .C(currBit[0]), 
         .D(currBit[3]), .Z(currPWMCountMax_15__N_230[12])) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i8724_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i3_4_lut (.A(\PWMArray[0][9] ), .B(currBit[0]), .C(currBit[3]), 
         .D(n12349), .Z(currPWMVal_15__N_213[0])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i3_4_lut.init = 16'h0800;
    LUT4 i1235_2_lut_3_lut_4_lut (.A(n12254), .B(n12241), .C(MATRIX_CURRROW[0]), 
         .D(n12281), .Z(n12[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(147[4] 185[11])
    defparam i1235_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1047_2_lut_3_lut_4_lut (.A(MATRIX_CURRROW[2]), .B(n12342), .C(MATRIX_CURRROW[4]), 
         .D(MATRIX_CURRROW[3]), .Z(currReadRow[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1047_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 mux_91_Mux_2_i3_4_lut (.A(\PWMArray[0][11] ), .B(n12337), .C(currBit[1]), 
         .D(currBit[0]), .Z(n3_adj_1219)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam mux_91_Mux_2_i3_4_lut.init = 16'hcac0;
    LUT4 i2_3_lut (.A(currBit[3]), .B(n6_adj_1240), .C(currBit[2]), .Z(currPWMVal_15__N_213[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i2_3_lut.init = 16'h4040;
    LUT4 currBit_0__bdd_4_lut (.A(currBit[0]), .B(currBit[3]), .C(\PWMArray[0][11] ), 
         .D(\PWMArray[0][12] ), .Z(n11718)) /* synthesis lut_function=(A (B (D))+!A !(B+!(C))) */ ;
    defparam currBit_0__bdd_4_lut.init = 16'h9810;
    PFUMX i8423 (.BLUT(n11312), .ALUT(n11313), .C0(currBit[1]), .Z(n11315));
    LUT4 mux_91_Mux_6_i6_3_lut (.A(n12336), .B(n12337), .C(currBit[1]), 
         .Z(n6_adj_1240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam mux_91_Mux_6_i6_3_lut.init = 16'hcaca;
    LUT4 i541_2_lut (.A(currBit[1]), .B(currBit[2]), .Z(n7_adj_1220)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(191[36:65])
    defparam i541_2_lut.init = 16'h6666;
    LUT4 MATRIX_ROWCLK_N_289_bdd_4_lut (.A(MATRIX_ROWCLK_N_289), .B(currPixel[0]), 
         .C(n12330), .D(currPixel[1]), .Z(n11924)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;
    defparam MATRIX_ROWCLK_N_289_bdd_4_lut.init = 16'h33c8;
    LUT4 n7302_bdd_3_lut (.A(currBit[2]), .B(currBit[0]), .C(currBit[1]), 
         .Z(n11724)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam n7302_bdd_3_lut.init = 16'h8181;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(currPixel[1]), .B(n12285), .C(currPixel[7]), 
         .D(n12275), .Z(n5345)) /* synthesis lut_function=(A (C)+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(157[10:27])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'he0a0;
    LUT4 i4684_2_lut (.A(currPWMCount_15__N_262[15]), .B(n12231), .Z(currPWMCount_15__N_149[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4684_2_lut.init = 16'h2222;
    LUT4 i4685_2_lut (.A(currPWMCount_15__N_262[14]), .B(n12231), .Z(currPWMCount_15__N_149[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4685_2_lut.init = 16'h2222;
    LUT4 i4686_2_lut (.A(currPWMCount_15__N_262[13]), .B(n12231), .Z(currPWMCount_15__N_149[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4686_2_lut.init = 16'h2222;
    LUT4 i4687_2_lut (.A(currPWMCount_15__N_262[12]), .B(n12231), .Z(currPWMCount_15__N_149[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4687_2_lut.init = 16'h2222;
    LUT4 i4688_2_lut (.A(currPWMCount_15__N_262[11]), .B(n12231), .Z(currPWMCount_15__N_149[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4688_2_lut.init = 16'h2222;
    CCU2D add_107_3 (.A0(currPWMCount[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9968), .COUT(n9969), .S0(currPWMCount_15__N_262[1]), 
          .S1(currPWMCount_15__N_262[2]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_3.INIT0 = 16'h5aaa;
    defparam add_107_3.INIT1 = 16'h5aaa;
    defparam add_107_3.INJECT1_0 = "NO";
    defparam add_107_3.INJECT1_1 = "NO";
    LUT4 i4689_2_lut (.A(currPWMCount_15__N_262[10]), .B(n12231), .Z(currPWMCount_15__N_149[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4689_2_lut.init = 16'h2222;
    LUT4 i8372_3_lut (.A(\BLUE[2] [6]), .B(\BLUE[2] [7]), .C(currBit[0]), 
         .Z(n11264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8372_3_lut.init = 16'hcaca;
    LUT4 i4696_2_lut (.A(currPWMCount_15__N_262[9]), .B(n12231), .Z(currPWMCount_15__N_149[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4696_2_lut.init = 16'h2222;
    LUT4 i8371_3_lut (.A(\BLUE[2] [4]), .B(\BLUE[2] [5]), .C(currBit[0]), 
         .Z(n11263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8371_3_lut.init = 16'hcaca;
    LUT4 i4697_2_lut (.A(currPWMCount_15__N_262[8]), .B(n12231), .Z(currPWMCount_15__N_149[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4697_2_lut.init = 16'h2222;
    LUT4 i6_2_lut (.A(currPWMCount[2]), .B(currPWMCount[7]), .Z(n22_adj_1222)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6_2_lut.init = 16'h8888;
    LUT4 i4698_2_lut (.A(currPWMCount_15__N_262[7]), .B(n12231), .Z(currPWMCount_15__N_149[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4698_2_lut.init = 16'h2222;
    LUT4 i4699_2_lut (.A(currPWMCount_15__N_262[6]), .B(n12231), .Z(currPWMCount_15__N_149[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4699_2_lut.init = 16'h2222;
    LUT4 i4567_2_lut (.A(currPWMCount_15__N_262[0]), .B(n12231), .Z(currPWMCount_15__N_149[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4567_2_lut.init = 16'h2222;
    LUT4 i8370_3_lut (.A(\BLUE[2] [2]), .B(\BLUE[2] [3]), .C(currBit[0]), 
         .Z(n11262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8370_3_lut.init = 16'hcaca;
    LUT4 i4700_2_lut (.A(currPWMCount_15__N_262[5]), .B(n12231), .Z(currPWMCount_15__N_149[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4700_2_lut.init = 16'h2222;
    LUT4 i8369_3_lut (.A(\BLUE[2] [0]), .B(\BLUE[2] [1]), .C(currBit[0]), 
         .Z(n11261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8369_3_lut.init = 16'hcaca;
    LUT4 i8365_3_lut (.A(\RED[3] [6]), .B(\RED[3] [7]), .C(currBit[0]), 
         .Z(n11257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8365_3_lut.init = 16'hcaca;
    LUT4 i8364_3_lut (.A(\RED[3] [4]), .B(\RED[3] [5]), .C(currBit[0]), 
         .Z(n11256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8364_3_lut.init = 16'hcaca;
    LUT4 i4701_2_lut (.A(currPWMCount_15__N_262[4]), .B(n12231), .Z(currPWMCount_15__N_149[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4701_2_lut.init = 16'h2222;
    LUT4 i4702_2_lut (.A(currPWMCount_15__N_262[3]), .B(n12231), .Z(currPWMCount_15__N_149[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4702_2_lut.init = 16'h2222;
    LUT4 i4703_2_lut (.A(currPWMCount_15__N_262[2]), .B(n12231), .Z(currPWMCount_15__N_149[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4703_2_lut.init = 16'h2222;
    LUT4 VRAM_READ_ADDR_7__I_0_189_2_lut_3_lut_4_lut (.A(currBit[0]), .B(n12349), 
         .C(VRAM_READ_ADDR[7]), .D(currBit[3]), .Z(VRAM_READ_ADDR_7__N_127)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam VRAM_READ_ADDR_7__I_0_189_2_lut_3_lut_4_lut.init = 16'h4bf0;
    LUT4 i4704_2_lut (.A(currPWMCount_15__N_262[1]), .B(n12231), .Z(currPWMCount_15__N_149[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(205[4] 209[11])
    defparam i4704_2_lut.init = 16'h2222;
    LUT4 i5_3_lut_rep_304 (.A(currPixel[3]), .B(n10_adj_1227), .C(currPixel[7]), 
         .Z(n12330)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i5_3_lut_rep_304.init = 16'hefef;
    PFUMX i8429 (.BLUT(n11317), .ALUT(n11318), .C0(currBit[1]), .Z(n11321));
    LUT4 i8363_3_lut (.A(\RED[3] [2]), .B(\RED[3] [3]), .C(currBit[0]), 
         .Z(n11255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8363_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_249_4_lut (.A(currPixel[3]), .B(n10_adj_1227), .C(currPixel[7]), 
         .D(currPixel[0]), .Z(n12275)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i1_2_lut_rep_249_4_lut.init = 16'hffef;
    LUT4 i2_3_lut_4_lut_adj_123 (.A(currPixel[3]), .B(n10_adj_1227), .C(currPixel[7]), 
         .D(n11924), .Z(PIXEL_CLOCK_enable_2)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i2_3_lut_4_lut_adj_123.init = 16'h1000;
    LUT4 i2717_2_lut_rep_209_3_lut_4_lut (.A(currPixel[7]), .B(n12249), 
         .C(n12281), .D(n12254), .Z(PIXEL_CLOCK_enable_24)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(147[4] 185[11])
    defparam i2717_2_lut_rep_209_3_lut_4_lut.init = 16'h8000;
    LUT4 i8362_3_lut (.A(\RED[3] [0]), .B(\RED[3] [1]), .C(currBit[0]), 
         .Z(n11254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8362_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_259_4_lut (.A(currPixel[3]), .B(n10_adj_1227), .C(currPixel[7]), 
         .D(currPixel[0]), .Z(n12285)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i1_2_lut_rep_259_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_124 (.A(currPixel[3]), .B(n10_adj_1227), 
         .C(currPixel[7]), .D(currPixel[0]), .Z(PIXEL_CLOCK_enable_3)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(177[10:27])
    defparam i1_2_lut_3_lut_4_lut_adj_124.init = 16'h1000;
    LUT4 i8358_3_lut (.A(\GREEN[3] [6]), .B(\GREEN[3] [7]), .C(currBit[0]), 
         .Z(n11250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8358_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_4_lut (.A(currPixel[7]), .B(currPixel[1]), .C(n10_adj_1227), 
         .D(currPixel[3]), .Z(PIXEL_CLOCK_enable_15)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i8357_3_lut (.A(\GREEN[3] [4]), .B(\GREEN[3] [5]), .C(currBit[0]), 
         .Z(n11249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8357_3_lut.init = 16'hcaca;
    LUT4 i8356_3_lut (.A(\GREEN[3] [2]), .B(\GREEN[3] [3]), .C(currBit[0]), 
         .Z(n11248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8356_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_125 (.A(currPixel[7]), .B(currPixel[1]), 
         .C(n12330), .D(currPixel[0]), .Z(PIXEL_CLOCK_enable_4)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(146[3] 186[10])
    defparam i1_2_lut_3_lut_4_lut_adj_125.init = 16'h0800;
    LUT4 i8355_3_lut (.A(\GREEN[3] [0]), .B(\GREEN[3] [1]), .C(currBit[0]), 
         .Z(n11247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8355_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_4_lut (.A(MATRIX_ROWCLK_N_289), .B(n12260), .C(n12249), 
         .D(currPixel[7]), .Z(PIXEL_CLOCK_enable_20)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(147[4] 185[11])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i8351_3_lut (.A(\BLUE[3] [6]), .B(\BLUE[3] [7]), .C(currBit[0]), 
         .Z(n11243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8351_3_lut.init = 16'hcaca;
    LUT4 i4652_2_lut_rep_307 (.A(currBit[0]), .B(currBit[1]), .Z(n12333)) /* synthesis lut_function=(A+(B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(191[36:65])
    defparam i4652_2_lut_rep_307.init = 16'heeee;
    LUT4 i1724_2_lut_3_lut (.A(currBit[0]), .B(currBit[1]), .C(currBit[2]), 
         .Z(n7_adj_1221)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(191[36:65])
    defparam i1724_2_lut_3_lut.init = 16'h1e1e;
    LUT4 mux_91_Mux_9_i8_3_lut_rep_308 (.A(\PWMArray[0][11] ), .B(\PWMArray[0][10] ), 
         .C(currBit[0]), .Z(n12334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam mux_91_Mux_9_i8_3_lut_rep_308.init = 16'hcaca;
    LUT4 i4872_2_lut_4_lut (.A(\PWMArray[0][11] ), .B(\PWMArray[0][10] ), 
         .C(currBit[0]), .D(n12349), .Z(n14_adj_1241)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i4872_2_lut_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_rep_309 (.A(currBit[0]), .B(\PWMArray[0][12] ), .Z(n12335)) /* synthesis lut_function=(A (B)) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i1_2_lut_rep_309.init = 16'h8888;
    LUT4 mux_91_Mux_10_i8_3_lut_rep_310 (.A(\PWMArray[0][12] ), .B(\PWMArray[0][11] ), 
         .C(currBit[0]), .Z(n12336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam mux_91_Mux_10_i8_3_lut_rep_310.init = 16'hcaca;
    LUT4 i1_2_lut_rep_280_4_lut (.A(\PWMArray[0][12] ), .B(\PWMArray[0][11] ), 
         .C(currBit[0]), .D(currBit[1]), .Z(n12306)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i1_2_lut_rep_280_4_lut.init = 16'hca00;
    LUT4 mux_91_Mux_8_i8_3_lut_rep_311 (.A(\PWMArray[0][10] ), .B(\PWMArray[0][9] ), 
         .C(currBit[0]), .Z(n12337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam mux_91_Mux_8_i8_3_lut_rep_311.init = 16'hcaca;
    LUT4 i4874_2_lut_4_lut (.A(\PWMArray[0][10] ), .B(\PWMArray[0][9] ), 
         .C(currBit[0]), .D(n12349), .Z(n14)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(190[28:57])
    defparam i4874_2_lut_4_lut.init = 16'hca00;
    LUT4 i9_4_lut (.A(currPWMCount[0]), .B(currPWMCount[1]), .C(currPWMCount[6]), 
         .D(currPWMCount[4]), .Z(n25)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    CCU2D add_107_15 (.A0(currPWMCount[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9974), .COUT(n9975), .S0(currPWMCount_15__N_262[13]), 
          .S1(currPWMCount_15__N_262[14]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_15.INIT0 = 16'h5aaa;
    defparam add_107_15.INIT1 = 16'h5aaa;
    defparam add_107_15.INJECT1_0 = "NO";
    defparam add_107_15.INJECT1_1 = "NO";
    LUT4 i7209_2_lut_3_lut (.A(currBit[1]), .B(currBit[0]), .C(currBit[2]), 
         .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i7209_2_lut_3_lut.init = 16'h7878;
    CCU2D add_107_13 (.A0(currPWMCount[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9973), .COUT(n9974), .S0(currPWMCount_15__N_262[11]), 
          .S1(currPWMCount_15__N_262[12]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_13.INIT0 = 16'h5aaa;
    defparam add_107_13.INIT1 = 16'h5aaa;
    defparam add_107_13.INJECT1_0 = "NO";
    defparam add_107_13.INJECT1_1 = "NO";
    LUT4 i7216_3_lut_4_lut (.A(currBit[1]), .B(currBit[0]), .C(currBit[2]), 
         .D(currBit[3]), .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i7216_3_lut_4_lut.init = 16'h7f80;
    LUT4 i8350_3_lut (.A(\BLUE[3] [4]), .B(\BLUE[3] [5]), .C(currBit[0]), 
         .Z(n11242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8350_3_lut.init = 16'hcaca;
    PFUMX i8430 (.BLUT(n11319), .ALUT(n11320), .C0(currBit[1]), .Z(n11322));
    LUT4 i1_2_lut_rep_223_3_lut (.A(currPixel[0]), .B(n12330), .C(currPixel[1]), 
         .Z(n12249)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam i1_2_lut_rep_223_3_lut.init = 16'hfefe;
    LUT4 i8349_3_lut (.A(\BLUE[3] [2]), .B(\BLUE[3] [3]), .C(currBit[0]), 
         .Z(n11241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8349_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_215_3_lut_4_lut (.A(currPixel[0]), .B(n12330), .C(currPixel[7]), 
         .D(currPixel[1]), .Z(n12241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam i1_2_lut_rep_215_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i7200_1_lut_rep_313 (.A(currBit[0]), .Z(n12339)) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i7200_1_lut_rep_313.init = 16'h5555;
    LUT4 i2_3_lut_4_lut_4_lut (.A(currBit[0]), .B(\PWMArray[0][12] ), .C(n12349), 
         .D(currBit[3]), .Z(currPWMVal_15__N_213[12])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_212_3_lut_4_lut_3_lut_4_lut (.A(currPixel[0]), .B(n12330), 
         .C(currPixel[7]), .D(currPixel[1]), .Z(PIXEL_CLOCK_enable_13)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam i1_2_lut_rep_212_3_lut_4_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i768_2_lut_rep_214_3_lut_4_lut (.A(currPixel[0]), .B(n12330), .C(currPixel[7]), 
         .D(currPixel[1]), .Z(n12240)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam i768_2_lut_rep_214_3_lut_4_lut.init = 16'h0010;
    LUT4 i4833_2_lut_rep_314 (.A(currBit[0]), .B(\PWMArray[0][9] ), .Z(n12340)) /* synthesis lut_function=(!(A+!(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i4833_2_lut_rep_314.init = 16'h4444;
    LUT4 i8629_2_lut_rep_228_3_lut (.A(currPixel[0]), .B(n12330), .C(currPixel[1]), 
         .Z(n12254)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(164[10:27])
    defparam i8629_2_lut_rep_228_3_lut.init = 16'h1010;
    CCU2D add_107_11 (.A0(currPWMCount[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(currPWMCount[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n9972), .COUT(n9973), .S0(currPWMCount_15__N_262[9]), 
          .S1(currPWMCount_15__N_262[10]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_11.INIT0 = 16'h5aaa;
    defparam add_107_11.INIT1 = 16'h5aaa;
    defparam add_107_11.INJECT1_0 = "NO";
    defparam add_107_11.INJECT1_1 = "NO";
    LUT4 mux_91_Mux_1_i3_4_lut_4_lut (.A(currBit[0]), .B(\PWMArray[0][9] ), 
         .C(currBit[1]), .D(\PWMArray[0][10] ), .Z(n3)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam mux_91_Mux_1_i3_4_lut_4_lut.init = 16'h4a40;
    PFUMX mux_91_Mux_7_i15 (.BLUT(n7_adj_1236), .ALUT(n14_adj_1237), .C0(currBit[3]), 
          .Z(currPWMVal_15__N_213[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;
    LUT4 i1028_2_lut_rep_316 (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .Z(n12342)) /* synthesis lut_function=(A (B)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1028_2_lut_rep_316.init = 16'h8888;
    LUT4 i1040_2_lut_3_lut_4_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[3]), .D(MATRIX_CURRROW[2]), .Z(currReadRow[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1040_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1035_2_lut_rep_285_3_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[2]), .Z(n12311)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1035_2_lut_rep_285_3_lut.init = 16'h8080;
    LUT4 i1042_2_lut_rep_258_3_lut_4_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[3]), .D(MATRIX_CURRROW[2]), .Z(n12284)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1042_2_lut_rep_258_3_lut_4_lut.init = 16'h8000;
    LUT4 i1033_2_lut_3_lut (.A(MATRIX_CURRROW[1]), .B(MATRIX_CURRROW[0]), 
         .C(MATRIX_CURRROW[2]), .Z(currReadRow[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam i1033_2_lut_3_lut.init = 16'h7878;
    LUT4 i8348_3_lut (.A(\BLUE[3] [0]), .B(\BLUE[3] [1]), .C(currBit[0]), 
         .Z(n11240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8348_3_lut.init = 16'hcaca;
    CCU2D add_107_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(currPWMCount[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n9968), .S1(currPWMCount_15__N_262[0]));   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/syn_arit.vhd(928[41:65])
    defparam add_107_1.INIT0 = 16'hF000;
    defparam add_107_1.INIT1 = 16'h5555;
    defparam add_107_1.INJECT1_0 = "NO";
    defparam add_107_1.INJECT1_1 = "NO";
    PFUMX mux_91_Mux_9_i15 (.BLUT(n7_adj_1235), .ALUT(n14_adj_1241), .C0(currBit[3]), 
          .Z(currPWMVal_15__N_213[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=6, LSE_RCOL=30, LSE_LLINE=139, LSE_RLINE=139 */ ;
    L6MUX21 i8354 (.D0(n11244), .D1(n11245), .SD(currBit[2]), .Z(n11246));
    L6MUX21 i8361 (.D0(n11251), .D1(n11252), .SD(currBit[2]), .Z(n11253));
    L6MUX21 i8368 (.D0(n11258), .D1(n11259), .SD(currBit[2]), .Z(n11260));
    LUT4 i10_4_lut (.A(currPWMCount[8]), .B(currPWMCount[3]), .C(currPWMCount[13]), 
         .D(currPWMCount[5]), .Z(n26)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i10_4_lut.init = 16'h8000;
    LUT4 n44_bdd_4_lut (.A(n37[1]), .B(n1095), .C(currPixel[1]), .D(n12275), 
         .Z(n12047)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A (((D)+!C)+!B))) */ ;
    defparam n44_bdd_4_lut.init = 16'h22e2;
    L6MUX21 i8375 (.D0(n11265), .D1(n11266), .SD(currBit[2]), .Z(n11267));
    L6MUX21 i8382 (.D0(n11272), .D1(n11273), .SD(currBit[2]), .Z(n11274));
    L6MUX21 i8389 (.D0(n11279), .D1(n11280), .SD(currBit[2]), .Z(n11281));
    Outputbuffer VRam (.VRAM_READ_ADDR_7__N_182(VRAM_WRITE_ADDR[7]), .\VRAM_ADDR[6] (\VRAM_ADDR[6] ), 
            .\VRAM_ADDR[5] (\VRAM_ADDR[5] ), .\VRAM_ADDR[4] (\VRAM_ADDR[4] ), 
            .\VRAM_ADDR[3] (\VRAM_ADDR[3] ), .\VRAM_ADDR[2] (\VRAM_ADDR[2] ), 
            .\VRAM_ADDR[1] (\VRAM_ADDR[1] ), .\VRAM_ADDR[0] (\VRAM_ADDR[0] ), 
            .\VRAM_READ_ADDR[7] (VRAM_READ_ADDR[7]), .\currPixel[6] (currPixel[6]), 
            .\currPixel[5] (currPixel[5]), .\currPixel[4] (currPixel[4]), 
            .\currPixel[3] (currPixel[3]), .\currPixel[2] (currPixel[2]), 
            .\currPixel[1] (currPixel[1]), .\currPixel[0] (currPixel[0]), 
            .n3028({n3028}), .n3027({n3027}), .VCC_net(VCC_net), .PIXEL_CLOCK_N_302(PIXEL_CLOCK_N_302), 
            .GND_net(GND_net), .VRAM_WC(VRAM_WC), .\BLUE[3] ({\BLUE[3] }), 
            .\GREEN[3] ({\GREEN[3] }), .n3035({n3035}), .n3034({n3034}), 
            .n3033({n3033}), .\RED[1] ({\RED[1] }), .\BLUE[0] ({\BLUE[0] }), 
            .\GREEN[0] ({\GREEN[0] }), .n3032({n3032}), .\RED[0] ({\RED[0] }), 
            .n3037({n3037}), .n3036({n3036}), .\BLUE[1] ({\BLUE[1] }), 
            .\GREEN[1] ({\GREEN[1] }), .n3030({n3030}), .n3029({n3029}), 
            .\GREEN[2] ({\GREEN[2] }), .\RED[2] ({\RED[2] }), .n3031({n3031}), 
            .\BLUE[2] ({\BLUE[2] }), .VRAM_DATA({VRAM_DATA}), .\RED[3] ({\RED[3] })) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    
endmodule
//
// Verilog Description of module Outputbuffer
//

module Outputbuffer (VRAM_READ_ADDR_7__N_182, \VRAM_ADDR[6] , \VRAM_ADDR[5] , 
            \VRAM_ADDR[4] , \VRAM_ADDR[3] , \VRAM_ADDR[2] , \VRAM_ADDR[1] , 
            \VRAM_ADDR[0] , \VRAM_READ_ADDR[7] , \currPixel[6] , \currPixel[5] , 
            \currPixel[4] , \currPixel[3] , \currPixel[2] , \currPixel[1] , 
            \currPixel[0] , n3028, n3027, VCC_net, PIXEL_CLOCK_N_302, 
            GND_net, VRAM_WC, \BLUE[3] , \GREEN[3] , n3035, n3034, 
            n3033, \RED[1] , \BLUE[0] , \GREEN[0] , n3032, \RED[0] , 
            n3037, n3036, \BLUE[1] , \GREEN[1] , n3030, n3029, \GREEN[2] , 
            \RED[2] , n3031, \BLUE[2] , VRAM_DATA, \RED[3] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input VRAM_READ_ADDR_7__N_182;
    input \VRAM_ADDR[6] ;
    input \VRAM_ADDR[5] ;
    input \VRAM_ADDR[4] ;
    input \VRAM_ADDR[3] ;
    input \VRAM_ADDR[2] ;
    input \VRAM_ADDR[1] ;
    input \VRAM_ADDR[0] ;
    input \VRAM_READ_ADDR[7] ;
    input \currPixel[6] ;
    input \currPixel[5] ;
    input \currPixel[4] ;
    input \currPixel[3] ;
    input \currPixel[2] ;
    input \currPixel[1] ;
    input \currPixel[0] ;
    input [9:0]n3028;
    input [9:0]n3027;
    input VCC_net;
    input PIXEL_CLOCK_N_302;
    input GND_net;
    input VRAM_WC;
    output [9:0]\BLUE[3] ;
    output [9:0]\GREEN[3] ;
    input [9:0]n3035;
    input [9:0]n3034;
    input [9:0]n3033;
    output [9:0]\RED[1] ;
    output [9:0]\BLUE[0] ;
    output [9:0]\GREEN[0] ;
    input [9:0]n3032;
    output [9:0]\RED[0] ;
    input [9:0]n3037;
    input [9:0]n3036;
    output [9:0]\BLUE[1] ;
    output [9:0]\GREEN[1] ;
    input [9:0]n3030;
    input [9:0]n3029;
    output [9:0]\GREEN[2] ;
    output [9:0]\RED[2] ;
    input [9:0]n3031;
    output [9:0]\BLUE[2] ;
    input [9:0]VRAM_DATA;
    output [9:0]\RED[3] ;
    
    wire PIXEL_CLOCK_N_302 /* synthesis is_inv_clock=1, is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(82[9:22])
    wire VRAM_WC /* synthesis is_clock=1 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/main.vhd(90[8:15])
    
    PDPW8KC Outputbuffer_0_6_0 (.DI0(n3027[8]), .DI1(n3027[9]), .DI2(n3028[0]), 
            .DI3(n3028[1]), .DI4(n3028[2]), .DI5(n3028[3]), .DI6(n3028[4]), 
            .DI7(n3028[5]), .DI8(n3028[6]), .DI9(n3028[7]), .DI10(n3028[8]), 
            .DI11(n3028[9]), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(\VRAM_ADDR[0] ), 
            .ADW1(\VRAM_ADDR[1] ), .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), 
            .ADW4(\VRAM_ADDR[4] ), .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), 
            .ADW7(VRAM_READ_ADDR_7__N_182), .ADW8(GND_net), .BE0(VCC_net), 
            .BE1(VCC_net), .CEW(VCC_net), .CLKW(VRAM_WC), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), 
            .ADR6(\currPixel[2] ), .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), 
            .ADR9(\currPixel[5] ), .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\BLUE[3] [7]), .DO1(\BLUE[3] [8]), .DO2(\BLUE[3] [9]), 
            .DO9(\GREEN[3] [8]), .DO10(\GREEN[3] [9]), .DO11(\BLUE[3] [0]), 
            .DO12(\BLUE[3] [1]), .DO13(\BLUE[3] [2]), .DO14(\BLUE[3] [3]), 
            .DO15(\BLUE[3] [4]), .DO16(\BLUE[3] [5]), .DO17(\BLUE[3] [6])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_6_0.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_6_0.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_6_0.REGMODE = "OUTREG";
    defparam Outputbuffer_0_6_0.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_6_0.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_6_0.GSR = "ENABLED";
    defparam Outputbuffer_0_6_0.RESETMODE = "SYNC";
    defparam Outputbuffer_0_6_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_6_0.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_6_0.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_6_0.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    PDPW8KC Outputbuffer_0_1_5 (.DI0(n3033[8]), .DI1(n3033[9]), .DI2(n3034[0]), 
            .DI3(n3034[1]), .DI4(n3034[2]), .DI5(n3034[3]), .DI6(n3034[4]), 
            .DI7(n3034[5]), .DI8(n3034[6]), .DI9(n3034[7]), .DI10(n3034[8]), 
            .DI11(n3034[9]), .DI12(n3035[0]), .DI13(n3035[1]), .DI14(n3035[2]), 
            .DI15(n3035[3]), .DI16(n3035[4]), .DI17(n3035[5]), .ADW0(\VRAM_ADDR[0] ), 
            .ADW1(\VRAM_ADDR[1] ), .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), 
            .ADW4(\VRAM_ADDR[4] ), .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), 
            .ADW7(VRAM_READ_ADDR_7__N_182), .ADW8(GND_net), .BE0(VCC_net), 
            .BE1(VCC_net), .CEW(VCC_net), .CLKW(VRAM_WC), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), 
            .ADR6(\currPixel[2] ), .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), 
            .ADR9(\currPixel[5] ), .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\BLUE[0] [7]), .DO1(\BLUE[0] [8]), .DO2(\BLUE[0] [9]), 
            .DO3(\RED[1] [0]), .DO4(\RED[1] [1]), .DO5(\RED[1] [2]), .DO6(\RED[1] [3]), 
            .DO7(\RED[1] [4]), .DO8(\RED[1] [5]), .DO9(\GREEN[0] [8]), 
            .DO10(\GREEN[0] [9]), .DO11(\BLUE[0] [0]), .DO12(\BLUE[0] [1]), 
            .DO13(\BLUE[0] [2]), .DO14(\BLUE[0] [3]), .DO15(\BLUE[0] [4]), 
            .DO16(\BLUE[0] [5]), .DO17(\BLUE[0] [6])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_1_5.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_1_5.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_1_5.REGMODE = "OUTREG";
    defparam Outputbuffer_0_1_5.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_1_5.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_1_5.GSR = "ENABLED";
    defparam Outputbuffer_0_1_5.RESETMODE = "SYNC";
    defparam Outputbuffer_0_1_5.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_1_5.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_1_5.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_1_5.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    PDPW8KC Outputbuffer_0_0_6 (.DI0(n3032[0]), .DI1(n3032[1]), .DI2(n3032[2]), 
            .DI3(n3032[3]), .DI4(n3032[4]), .DI5(n3032[5]), .DI6(n3032[6]), 
            .DI7(n3032[7]), .DI8(n3032[8]), .DI9(n3032[9]), .DI10(n3033[0]), 
            .DI11(n3033[1]), .DI12(n3033[2]), .DI13(n3033[3]), .DI14(n3033[4]), 
            .DI15(n3033[5]), .DI16(n3033[6]), .DI17(n3033[7]), .ADW0(\VRAM_ADDR[0] ), 
            .ADW1(\VRAM_ADDR[1] ), .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), 
            .ADW4(\VRAM_ADDR[4] ), .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), 
            .ADW7(VRAM_READ_ADDR_7__N_182), .ADW8(GND_net), .BE0(VCC_net), 
            .BE1(VCC_net), .CEW(VCC_net), .CLKW(VRAM_WC), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), 
            .ADR6(\currPixel[2] ), .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), 
            .ADR9(\currPixel[5] ), .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\RED[0] [9]), .DO1(\GREEN[0] [0]), .DO2(\GREEN[0] [1]), 
            .DO3(\GREEN[0] [2]), .DO4(\GREEN[0] [3]), .DO5(\GREEN[0] [4]), 
            .DO6(\GREEN[0] [5]), .DO7(\GREEN[0] [6]), .DO8(\GREEN[0] [7]), 
            .DO9(\RED[0] [0]), .DO10(\RED[0] [1]), .DO11(\RED[0] [2]), 
            .DO12(\RED[0] [3]), .DO13(\RED[0] [4]), .DO14(\RED[0] [5]), 
            .DO15(\RED[0] [6]), .DO16(\RED[0] [7]), .DO17(\RED[0] [8])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_0_6.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_0_6.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_0_6.REGMODE = "OUTREG";
    defparam Outputbuffer_0_0_6.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_0_6.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_0_6.GSR = "ENABLED";
    defparam Outputbuffer_0_0_6.RESETMODE = "SYNC";
    defparam Outputbuffer_0_0_6.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_0_6.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_0_6.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_0_6.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    PDPW8KC Outputbuffer_0_2_4 (.DI0(n3035[6]), .DI1(n3035[7]), .DI2(n3035[8]), 
            .DI3(n3035[9]), .DI4(n3036[0]), .DI5(n3036[1]), .DI6(n3036[2]), 
            .DI7(n3036[3]), .DI8(n3036[4]), .DI9(n3036[5]), .DI10(n3036[6]), 
            .DI11(n3036[7]), .DI12(n3036[8]), .DI13(n3036[9]), .DI14(n3037[0]), 
            .DI15(n3037[1]), .DI16(n3037[2]), .DI17(n3037[3]), .ADW0(\VRAM_ADDR[0] ), 
            .ADW1(\VRAM_ADDR[1] ), .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), 
            .ADW4(\VRAM_ADDR[4] ), .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), 
            .ADW7(VRAM_READ_ADDR_7__N_182), .ADW8(GND_net), .BE0(VCC_net), 
            .BE1(VCC_net), .CEW(VCC_net), .CLKW(VRAM_WC), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), 
            .ADR6(\currPixel[2] ), .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), 
            .ADR9(\currPixel[5] ), .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\GREEN[1] [5]), .DO1(\GREEN[1] [6]), .DO2(\GREEN[1] [7]), 
            .DO3(\GREEN[1] [8]), .DO4(\GREEN[1] [9]), .DO5(\BLUE[1] [0]), 
            .DO6(\BLUE[1] [1]), .DO7(\BLUE[1] [2]), .DO8(\BLUE[1] [3]), 
            .DO9(\RED[1] [6]), .DO10(\RED[1] [7]), .DO11(\RED[1] [8]), 
            .DO12(\RED[1] [9]), .DO13(\GREEN[1] [0]), .DO14(\GREEN[1] [1]), 
            .DO15(\GREEN[1] [2]), .DO16(\GREEN[1] [3]), .DO17(\GREEN[1] [4])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_2_4.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_2_4.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_2_4.REGMODE = "OUTREG";
    defparam Outputbuffer_0_2_4.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_2_4.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_2_4.GSR = "ENABLED";
    defparam Outputbuffer_0_2_4.RESETMODE = "SYNC";
    defparam Outputbuffer_0_2_4.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_2_4.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_2_4.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_2_4.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    PDPW8KC Outputbuffer_0_3_3 (.DI0(n3037[4]), .DI1(n3037[5]), .DI2(n3037[6]), 
            .DI3(n3037[7]), .DI4(n3037[8]), .DI5(n3037[9]), .DI6(n3029[0]), 
            .DI7(n3029[1]), .DI8(n3029[2]), .DI9(n3029[3]), .DI10(n3029[4]), 
            .DI11(n3029[5]), .DI12(n3029[6]), .DI13(n3029[7]), .DI14(n3029[8]), 
            .DI15(n3029[9]), .DI16(n3030[0]), .DI17(n3030[1]), .ADW0(\VRAM_ADDR[0] ), 
            .ADW1(\VRAM_ADDR[1] ), .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), 
            .ADW4(\VRAM_ADDR[4] ), .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), 
            .ADW7(VRAM_READ_ADDR_7__N_182), .ADW8(GND_net), .BE0(VCC_net), 
            .BE1(VCC_net), .CEW(VCC_net), .CLKW(VRAM_WC), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), 
            .ADR6(\currPixel[2] ), .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), 
            .ADR9(\currPixel[5] ), .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\RED[2] [3]), .DO1(\RED[2] [4]), .DO2(\RED[2] [5]), .DO3(\RED[2] [6]), 
            .DO4(\RED[2] [7]), .DO5(\RED[2] [8]), .DO6(\RED[2] [9]), .DO7(\GREEN[2] [0]), 
            .DO8(\GREEN[2] [1]), .DO9(\BLUE[1] [4]), .DO10(\BLUE[1] [5]), 
            .DO11(\BLUE[1] [6]), .DO12(\BLUE[1] [7]), .DO13(\BLUE[1] [8]), 
            .DO14(\BLUE[1] [9]), .DO15(\RED[2] [0]), .DO16(\RED[2] [1]), 
            .DO17(\RED[2] [2])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_3_3.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_3_3.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_3_3.REGMODE = "OUTREG";
    defparam Outputbuffer_0_3_3.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_3_3.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_3_3.GSR = "ENABLED";
    defparam Outputbuffer_0_3_3.RESETMODE = "SYNC";
    defparam Outputbuffer_0_3_3.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_3_3.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_3_3.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_3_3.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    PDPW8KC Outputbuffer_0_4_2 (.DI0(n3030[2]), .DI1(n3030[3]), .DI2(n3030[4]), 
            .DI3(n3030[5]), .DI4(n3030[6]), .DI5(n3030[7]), .DI6(n3030[8]), 
            .DI7(n3030[9]), .DI8(n3031[0]), .DI9(n3031[1]), .DI10(n3031[2]), 
            .DI11(n3031[3]), .DI12(n3031[4]), .DI13(n3031[5]), .DI14(n3031[6]), 
            .DI15(n3031[7]), .DI16(n3031[8]), .DI17(n3031[9]), .ADW0(\VRAM_ADDR[0] ), 
            .ADW1(\VRAM_ADDR[1] ), .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), 
            .ADW4(\VRAM_ADDR[4] ), .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), 
            .ADW7(VRAM_READ_ADDR_7__N_182), .ADW8(GND_net), .BE0(VCC_net), 
            .BE1(VCC_net), .CEW(VCC_net), .CLKW(VRAM_WC), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), 
            .ADR6(\currPixel[2] ), .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), 
            .ADR9(\currPixel[5] ), .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\BLUE[2] [1]), .DO1(\BLUE[2] [2]), .DO2(\BLUE[2] [3]), 
            .DO3(\BLUE[2] [4]), .DO4(\BLUE[2] [5]), .DO5(\BLUE[2] [6]), 
            .DO6(\BLUE[2] [7]), .DO7(\BLUE[2] [8]), .DO8(\BLUE[2] [9]), 
            .DO9(\GREEN[2] [2]), .DO10(\GREEN[2] [3]), .DO11(\GREEN[2] [4]), 
            .DO12(\GREEN[2] [5]), .DO13(\GREEN[2] [6]), .DO14(\GREEN[2] [7]), 
            .DO15(\GREEN[2] [8]), .DO16(\GREEN[2] [9]), .DO17(\BLUE[2] [0])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_4_2.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_4_2.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_4_2.REGMODE = "OUTREG";
    defparam Outputbuffer_0_4_2.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_4_2.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_4_2.GSR = "ENABLED";
    defparam Outputbuffer_0_4_2.RESETMODE = "SYNC";
    defparam Outputbuffer_0_4_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_4_2.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_4_2.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_4_2.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    PDPW8KC Outputbuffer_0_5_1 (.DI0(VRAM_DATA[0]), .DI1(VRAM_DATA[1]), 
            .DI2(VRAM_DATA[2]), .DI3(VRAM_DATA[3]), .DI4(VRAM_DATA[4]), 
            .DI5(VRAM_DATA[5]), .DI6(VRAM_DATA[6]), .DI7(VRAM_DATA[7]), 
            .DI8(VRAM_DATA[8]), .DI9(VRAM_DATA[9]), .DI10(n3027[0]), .DI11(n3027[1]), 
            .DI12(n3027[2]), .DI13(n3027[3]), .DI14(n3027[4]), .DI15(n3027[5]), 
            .DI16(n3027[6]), .DI17(n3027[7]), .ADW0(\VRAM_ADDR[0] ), .ADW1(\VRAM_ADDR[1] ), 
            .ADW2(\VRAM_ADDR[2] ), .ADW3(\VRAM_ADDR[3] ), .ADW4(\VRAM_ADDR[4] ), 
            .ADW5(\VRAM_ADDR[5] ), .ADW6(\VRAM_ADDR[6] ), .ADW7(VRAM_READ_ADDR_7__N_182), 
            .ADW8(GND_net), .BE0(VCC_net), .BE1(VCC_net), .CEW(VCC_net), 
            .CLKW(VRAM_WC), .CSW0(VCC_net), .CSW1(GND_net), .CSW2(GND_net), 
            .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), .ADR3(GND_net), 
            .ADR4(\currPixel[0] ), .ADR5(\currPixel[1] ), .ADR6(\currPixel[2] ), 
            .ADR7(\currPixel[3] ), .ADR8(\currPixel[4] ), .ADR9(\currPixel[5] ), 
            .ADR10(\currPixel[6] ), .ADR11(\VRAM_READ_ADDR[7] ), .ADR12(GND_net), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(PIXEL_CLOCK_N_302), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(\RED[3] [9]), 
            .DO1(\GREEN[3] [0]), .DO2(\GREEN[3] [1]), .DO3(\GREEN[3] [2]), 
            .DO4(\GREEN[3] [3]), .DO5(\GREEN[3] [4]), .DO6(\GREEN[3] [5]), 
            .DO7(\GREEN[3] [6]), .DO8(\GREEN[3] [7]), .DO9(\RED[3] [0]), 
            .DO10(\RED[3] [1]), .DO11(\RED[3] [2]), .DO12(\RED[3] [3]), 
            .DO13(\RED[3] [4]), .DO14(\RED[3] [5]), .DO15(\RED[3] [6]), 
            .DO16(\RED[3] [7]), .DO17(\RED[3] [8])) /* synthesis MEM_LPC_FILE="Outputbuffer.lpc", MEM_INIT_FILE="INIT_ALL_1s", syn_instantiated=1, LSE_LINE_FILE_ID=22, LSE_LCOL=8, LSE_RCOL=20, LSE_LLINE=246, LSE_RLINE=246 */ ;   // d:/onedrive/lattice diamond projects/wallpanel_fpga/matrixdriver.vhd(246[8:20])
    defparam Outputbuffer_0_5_1.DATA_WIDTH_W = 18;
    defparam Outputbuffer_0_5_1.DATA_WIDTH_R = 18;
    defparam Outputbuffer_0_5_1.REGMODE = "OUTREG";
    defparam Outputbuffer_0_5_1.CSDECODE_W = "0b001";
    defparam Outputbuffer_0_5_1.CSDECODE_R = "0b000";
    defparam Outputbuffer_0_5_1.GSR = "ENABLED";
    defparam Outputbuffer_0_5_1.RESETMODE = "SYNC";
    defparam Outputbuffer_0_5_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam Outputbuffer_0_5_1.INIT_DATA = "STATIC";
    defparam Outputbuffer_0_5_1.INITVAL_00 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_01 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_02 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_03 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_04 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_05 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_06 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_07 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_08 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_09 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_0A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_0B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_0C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_0D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_0E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_0F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_10 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_11 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_12 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_13 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_14 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_15 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_16 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_17 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_18 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_19 = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_1A = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_1B = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_1C = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_1D = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_1E = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    defparam Outputbuffer_0_5_1.INITVAL_1F = "0xFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    
endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Sun Jan 10 17:32:53 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Sun Jan 10 17:32:52 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Sun Jan 10 17:49:31 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Sun Jan 10 17:49:30 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Sun Jan 10 18:07:24 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Sun Jan 10 18:07:23 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 14:04:04 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 14:04:03 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 14:07:22 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 14:07:21 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 14:10:46 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 14:10:45 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 14:22:54 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 14:22:53 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 14:56:09 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 14:56:08 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 15:01:18 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 15:01:17 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 15:56:05 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 15:56:04 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 16:00:24 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 16:00:23 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 16:04:14 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 16:04:13 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 3.9 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type sdpram -num_rows 32 -data_width 2 -pipe_final_output -memformat bin -n pmi_distributed_dpramXbnoner25328de3a5d -pmi -lang verilog  */
/* Mon Jan 11 16:08:04 2021 */


`timescale 1 ns / 1 ps
module pmi_distributed_dpramXbnoner25328de3a5d (WrAddress, Data, WrClock, 
    WE, WrClockEn, RdAddress, RdClock, RdClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [1:0] Data;
    input wire WrClock;
    input wire WE;
    input wire WrClockEn;
    input wire [4:0] RdAddress;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    output wire [1:0] Q;

    wire waddr4_inv;
    wire dataout1_ffin;
    wire dataout0_ffin;
    wire mdL0_0_1;
    wire mdL0_0_0;
    wire dec0_wre3;
    wire mdL0_1_1;
    wire mdL0_1_0;
    wire dec1_wre7;
    wire scuba_vhi;

    INV INV_0 (.A(WrAddress[4]), .Z(waddr4_inv));

    defparam LUT4_1.initval =  16'h8000 ;
    ROM16X1A LUT4_1 (.AD3(WE), .AD2(WrClockEn), .AD1(waddr4_inv), .AD0(scuba_vhi), 
        .DO0(dec0_wre3));

    defparam LUT4_0.initval =  16'h8000 ;
    ROM16X1A LUT4_0 (.AD3(WE), .AD2(WrClockEn), .AD1(WrAddress[4]), .AD0(scuba_vhi), 
        .DO0(dec1_wre7));

    FD1P3DX FF_1 (.D(dataout1_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[1]))
             /* synthesis GSR="ENABLED" */;

    FD1P3DX FF_0 (.D(dataout0_ffin), .SP(RdClockEn), .CK(RdClock), .CD(Reset), 
        .Q(Q[0]))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_1 (.D0(mdL0_0_1), .D1(mdL0_1_1), .SD(RdAddress[4]), .Z(dataout1_ffin));

    MUX21 mux_0 (.D0(mdL0_0_0), .D1(mdL0_1_0), .SD(RdAddress[4]), .Z(dataout0_ffin));

    defparam mem_0_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_0_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec0_wre3), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_0_0), .DO1(mdL0_0_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(0-15)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_0_0" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam mem_1_0.initval = "0x0000000000000000" ;
    DPR16X4C mem_1_0 (.DI0(Data[0]), .DI1(Data[1]), .DI2(scuba_vhi), .DI3(scuba_vhi), 
        .WCK(WrClock), .WRE(dec1_wre7), .RAD0(RdAddress[0]), .RAD1(RdAddress[1]), 
        .RAD2(RdAddress[2]), .RAD3(RdAddress[3]), .WAD0(WrAddress[0]), .WAD1(WrAddress[1]), 
        .WAD2(WrAddress[2]), .WAD3(WrAddress[3]), .DO0(mdL0_1_0), .DO1(mdL0_1_1), 
        .DO2(), .DO3())
             /* synthesis MEM_INIT_FILE="(16-31)(0-1)" */
             /* synthesis MEM_LPC_FILE="pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B" */
             /* synthesis COMP="mem_1_0" */;



    // exemplar begin
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar attribute mem_0_0 MEM_INIT_FILE (0-15)(0-1)
    // exemplar attribute mem_0_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_0_0 COMP mem_0_0
    // exemplar attribute mem_1_0 MEM_INIT_FILE (16-31)(0-1)
    // exemplar attribute mem_1_0 MEM_LPC_FILE pmi_distributed_dpramXbnoner25328de3a5d__PMI__32__2__2B
    // exemplar attribute mem_1_0 COMP mem_1_0
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.11.0.396.4 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.11_x64/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo3c00f -type bram -wp 10 -rp 0011 -data_width 146 -num_rows 1024 -rdata_width 146 -read_reg1 outreg -gsr DISABLED -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr146101024146101024123cc668 -pmi -lang verilog  */
/* Mon Jan 11 16:08:03 2021 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr146101024146101024123cc668 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] WrAddress;
    input wire [9:0] RdAddress;
    input wire [145:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [145:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[8]), .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), 
        .DOB3(Q[3]), .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[17]), .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), 
        .DOB4(Q[13]), .DOB3(Q[12]), .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[26]), .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), 
        .DOB4(Q[22]), .DOB3(Q[21]), .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[35]), .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), 
        .DOB4(Q[31]), .DOB3(Q[30]), .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[44]), .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), 
        .DOB4(Q[40]), .DOB3(Q[39]), .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[53]), .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), 
        .DOB4(Q[49]), .DOB3(Q[48]), .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[62]), .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), 
        .DOB4(Q[58]), .DOB3(Q[57]), .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[71]), .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), 
        .DOB4(Q[67]), .DOB3(Q[66]), .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[80]), .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), 
        .DOB4(Q[76]), .DOB3(Q[75]), .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[89]), .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), 
        .DOB4(Q[85]), .DOB3(Q[84]), .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 (.DIA8(Data[98]), 
        .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), .DIA4(Data[94]), 
        .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[98]), .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), 
        .DOB4(Q[94]), .DOB3(Q[93]), .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 (.DIA8(Data[107]), 
        .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), .DIA4(Data[103]), 
        .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), .DIA0(Data[99]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[107]), .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), 
        .DOB4(Q[103]), .DOB3(Q[102]), .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 (.DIA8(Data[116]), 
        .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), .DIA4(Data[112]), 
        .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), .DIA0(Data[108]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[116]), .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), 
        .DOB4(Q[112]), .DOB3(Q[111]), .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 (.DIA8(Data[125]), 
        .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), .DIA4(Data[121]), 
        .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), .DIA0(Data[117]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[125]), .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), 
        .DOB4(Q[121]), .DOB3(Q[120]), .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 (.DIA8(Data[134]), 
        .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), .DIA4(Data[130]), 
        .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), .DIA0(Data[126]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[134]), .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), 
        .DOB4(Q[130]), .DOB3(Q[129]), .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 (.DIA8(Data[143]), 
        .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), .DIA4(Data[139]), 
        .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), .DIA0(Data[135]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(Q[143]), .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), 
        .DOB4(Q[139]), .DOB3(Q[138]), .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[145]), .DIA0(Data[144]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(scuba_vlo), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr146101024146101024123cc668__PMIP__1024__146__146B
    // exemplar attribute pmi_ram_dpXbnonesadr146101024146101024123cc668_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
